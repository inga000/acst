.suckt  symmetrical_op_amp89 ibias in1 in2 out sourceNmos sourcePmos
mSymmetricalFirstStageLoad1 out2FirstStage out2FirstStage out1FirstStage out1FirstStage nmos
mSymmetricalFirstStageLoad2 out1FirstStage out1FirstStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageLoad3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage nmos
mSymmetricalFirstStageLoad4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSymmetricalFirstStageTransconductor6 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSymmetricalFirstStageTransconductor7 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1Transconductor8 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mSecondStage1Transconductor9 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias10 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mSecondStage1StageBias11 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias12 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias13 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mMainBias16 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp89

