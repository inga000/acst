** Name: two_stage_single_output_op_amp_203_8

.MACRO two_stage_single_output_op_amp_203_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=17e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
m3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=16e-6
m5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
m6 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=221e-6
m7 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=16e-6
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=104e-6
m9 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=114e-6
m10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=115e-6
m11 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
m12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=104e-6
m13 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=47e-6
m14 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
m15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=522e-6
m16 outFirstStage outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=50e-6
m17 FirstStageYout1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=50e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10.8001e-12
.EOM two_stage_single_output_op_amp_203_8

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 3.56701 mW
** Area: 8538 (mu_m)^2
** Transit frequency: 4.30901 MHz
** Transit frequency with error factor: 4.28027 MHz
** Slew rate: 4.06069 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.84001 V
** VoutMin: 0.800001 V
** VcmMax: 4.71001 V
** VcmMin: 1.35001 V


** Expected Currents: 
** NormalTransistorNmos: 4.37181e+07 muA
** DiodeTransistorNmos: 1.92359e+08 muA
** NormalTransistorNmos: 1.9236e+08 muA
** NormalTransistorNmos: 1.92359e+08 muA
** DiodeTransistorNmos: 1.9236e+08 muA
** NormalTransistorPmos: -2.14368e+08 muA
** NormalTransistorPmos: -2.14368e+08 muA
** NormalTransistorNmos: 4.40191e+07 muA
** NormalTransistorNmos: 4.40181e+07 muA
** NormalTransistorNmos: 2.20101e+07 muA
** NormalTransistorNmos: 2.20101e+07 muA
** NormalTransistorNmos: 2.30865e+08 muA
** NormalTransistorNmos: 2.30864e+08 muA
** NormalTransistorPmos: -2.30864e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -4.37189e+07 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.27801  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 3.74001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.06101  V
** innerStageBias: 0.505001  V
** innerTransistorStack1Load1: 1.06101  V
** out1: 2.21601  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.492001  V


.END