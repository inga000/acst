** Name: two_stage_single_output_op_amp_76_7

.MACRO two_stage_single_output_op_amp_76_7 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
m2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=71e-6
m3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=13e-6
m4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=52e-6
m5 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=56e-6
m6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=38e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=24e-6
m8 out inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=198e-6
m9 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=94e-6
m10 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=56e-6
m11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=16e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=16e-6
m13 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=52e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=13e-6
m15 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=70e-6
m16 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=521e-6
m17 out outFirstStage sourcePmos sourcePmos pmos4 L=10e-6 W=562e-6
m18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=67e-6
m19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=14e-6
m20 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=67e-6
m21 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=83e-6
m22 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=83e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 5e-12
.EOM two_stage_single_output_op_amp_76_7

** Expected Performance Values: 
** Gain: 112 dB
** Power consumption: 4.56201 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 2.65001 MHz
** Transit frequency with error factor: 2.64998 MHz
** Slew rate: 4.64073 V/mu_s
** Phase margin: 60.1606°
** CMRR: 136 dB
** VoutMax: 4.25 V
** VoutMin: 0.590001 V
** VcmMax: 5.10001 V
** VcmMin: 1.42001 V


** Expected Currents: 
** NormalTransistorPmos: -5.90799e+06 muA
** NormalTransistorPmos: -2.16329e+08 muA
** NormalTransistorPmos: -2.93629e+07 muA
** NormalTransistorPmos: -2.33809e+07 muA
** NormalTransistorPmos: -3.50709e+07 muA
** NormalTransistorPmos: -2.33809e+07 muA
** NormalTransistorPmos: -3.50709e+07 muA
** DiodeTransistorNmos: 2.33801e+07 muA
** NormalTransistorNmos: 2.33801e+07 muA
** NormalTransistorNmos: 2.33801e+07 muA
** NormalTransistorNmos: 2.33811e+07 muA
** DiodeTransistorNmos: 2.33801e+07 muA
** NormalTransistorNmos: 1.16911e+07 muA
** NormalTransistorNmos: 1.16911e+07 muA
** NormalTransistorNmos: 5.70621e+08 muA
** NormalTransistorPmos: -5.7062e+08 muA
** DiodeTransistorNmos: 5.90701e+06 muA
** NormalTransistorNmos: 5.90601e+06 muA
** DiodeTransistorNmos: 2.1633e+08 muA
** DiodeTransistorNmos: 2.93621e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.977001  V
** inputVoltageBiasXXnXX3: 0.991001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.13601  V
** outSourceVoltageBiasXXnXX1: 0.568001  V
** outSourceVoltageBiasXXpXX1: 4.13001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.410001  V
** out1: 0.615001  V
** sourceGCC1: 4.16601  V
** sourceGCC2: 4.16601  V
** sourceTransconductance: 1.81501  V
** inner: 0.567001  V


.END