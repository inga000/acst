** Name: one_stage_single_output_op_amp45

.MACRO one_stage_single_output_op_amp45 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=5e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=163e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=79e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=115e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=115e-6
mMainBias9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=195e-6
mMainBias10 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=60e-6
mFoldedCascodeFirstStageLoad11 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=163e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=157e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=157e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=113e-6
mFoldedCascodeFirstStageLoad16 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=25e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp45

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 2.44301 mW
** Area: 3966 (mu_m)^2
** Transit frequency: 2.75401 MHz
** Transit frequency with error factor: 2.7539 MHz
** Slew rate: 3.50001 V/mu_s
** Phase margin: 89.3815°
** CMRR: 140 dB
** VoutMax: 4.45001 V
** VoutMin: 0.75 V
** VcmMax: 3.68001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.92914e+08 muA
** NormalTransistorNmos: 6.00471e+07 muA
** NormalTransistorNmos: 7.00581e+07 muA
** NormalTransistorNmos: 1.12815e+08 muA
** NormalTransistorNmos: 7.00551e+07 muA
** NormalTransistorNmos: 1.12814e+08 muA
** DiodeTransistorPmos: -7.00569e+07 muA
** NormalTransistorPmos: -7.00559e+07 muA
** NormalTransistorPmos: -7.00569e+07 muA
** NormalTransistorPmos: -8.55149e+07 muA
** NormalTransistorPmos: -4.27569e+07 muA
** NormalTransistorPmos: -4.27569e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.92913e+08 muA
** DiodeTransistorPmos: -6.00479e+07 muA


** Expected Voltages: 
** ibias: 1.18001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** inputVoltageBiasXXpXX2: 3.93001  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.64501  V
** out1: 4.28101  V
** sourceGCC1: 0.587001  V
** sourceGCC2: 0.587001  V
** sourceTransconductance: 3.31001  V


.END