** Name: two_stage_single_output_op_amp_9_11

.MACRO two_stage_single_output_op_amp_9_11 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=78e-6
m3 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=240e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=71e-6
m5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=333e-6
m6 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=6e-6 W=133e-6
m7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=11e-6
m8 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=300e-6
m9 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=325e-6
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=11e-6
m11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=131e-6
m12 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=574e-6
m13 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=591e-6
m14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=213e-6
m15 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=440e-6
m16 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=333e-6
m17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=221e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 15.2001e-12
.EOM two_stage_single_output_op_amp_9_11

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 10.4431 mW
** Area: 11357 (mu_m)^2
** Transit frequency: 3.81701 MHz
** Transit frequency with error factor: 3.81207 MHz
** Slew rate: 9.43341 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 101 dB
** posPSRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 0.740001 V
** VcmMax: 4.46001 V
** VcmMin: 0.960001 V


** Expected Currents: 
** NormalTransistorNmos: 3.34128e+08 muA
** NormalTransistorNmos: 3.60445e+08 muA
** NormalTransistorPmos: -6.01488e+08 muA
** NormalTransistorPmos: -7.20369e+07 muA
** NormalTransistorPmos: -7.20369e+07 muA
** DiodeTransistorPmos: -7.20369e+07 muA
** NormalTransistorNmos: 1.44073e+08 muA
** NormalTransistorNmos: 7.20361e+07 muA
** NormalTransistorNmos: 7.20361e+07 muA
** NormalTransistorNmos: 6.38556e+08 muA
** NormalTransistorNmos: 6.38555e+08 muA
** NormalTransistorPmos: -6.38555e+08 muA
** NormalTransistorPmos: -6.38556e+08 muA
** DiodeTransistorNmos: 6.01489e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.34127e+08 muA
** DiodeTransistorPmos: -3.60444e+08 muA


** Expected Voltages: 
** ibias: 0.567001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.03201  V
** outVoltageBiasXXnXX1: 1.14801  V
** outVoltageBiasXXpXX0: 3.81501  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.24501  V
** out1: 3.48601  V
** sourceTransconductance: 1.70001  V
** innerStageBias: 0.162001  V
** innerTransconductance: 4.59601  V


.END