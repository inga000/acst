** Name: two_stage_single_output_op_amp_205_7

.MACRO two_stage_single_output_op_amp_205_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=10e-6 W=52e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=16e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=19e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=35e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=10e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=60e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=485e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=10e-6 W=52e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=35e-6
mSimpleFirstStageLoad14 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=292e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=194e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=194e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=262e-6
mSimpleFirstStageLoad18 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=292e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=125e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.5e-12
.EOM two_stage_single_output_op_amp_205_7

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 9.51301 mW
** Area: 7147 (mu_m)^2
** Transit frequency: 4.28201 MHz
** Transit frequency with error factor: 4.28033 MHz
** Slew rate: 4.03578 V/mu_s
** Phase margin: 60.1606°
** CMRR: 119 dB
** VoutMax: 4.25 V
** VoutMin: 0.400001 V
** VcmMax: 4.98001 V
** VcmMin: 1.54001 V


** Expected Currents: 
** NormalTransistorPmos: -1.26733e+08 muA
** NormalTransistorPmos: -5.04509e+07 muA
** DiodeTransistorNmos: 1.82439e+08 muA
** NormalTransistorNmos: 1.8244e+08 muA
** NormalTransistorNmos: 1.8244e+08 muA
** DiodeTransistorNmos: 1.8244e+08 muA
** NormalTransistorPmos: -1.95771e+08 muA
** NormalTransistorPmos: -1.95772e+08 muA
** NormalTransistorPmos: -1.95772e+08 muA
** NormalTransistorPmos: -1.95772e+08 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 2.66641e+07 muA
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 1.31381e+09 muA
** NormalTransistorPmos: -1.3138e+09 muA
** DiodeTransistorNmos: 1.26734e+08 muA
** DiodeTransistorNmos: 5.04501e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.15101  V
** outVoltageBiasXXnXX2: 0.803001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.10401  V
** innerStageBias: 0.568001  V
** innerTransistorStack1Load1: 1.05301  V
** innerTransistorStack1Load2: 4.15501  V
** innerTransistorStack2Load1: 1.05201  V
** innerTransistorStack2Load2: 4.15501  V
** sourceTransconductance: 1.94501  V


.END