.suckt  two_stage_fully_differential_op_amp_12_11 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_3 inputVoltageBiasXXpXX3 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_4 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_5 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_Load_6 outFeedback outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m_FullyDifferential_FeedbackdStage_StageBias_8 FeedbackStageYinnerStageBias1 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m_FullyDifferential_FeedbackdStage_StageBias_10 FeedbackStageYinnerStageBias2 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackStage_Transconductor_11 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FeedbackStage_Transconductor_14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FirstStage_Load_15 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m_FullyDifferential_FirstStage_Load_16 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m_FullyDifferential_FirstStage_Load_17 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m_FullyDifferential_FirstStage_Load_18 FirstStageYinnerTransistorStack1Load2 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_19 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m_FullyDifferential_FirstStage_Load_20 FirstStageYinnerTransistorStack2Load2 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_StageBias_21 sourceTransconductance inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Transconductor_22 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m_FullyDifferential_FirstStage_Transconductor_23 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_StageBias_24 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias nmos
m_FullyDifferential_SecondStage1_StageBias_25 SecondStage1YinnerStageBias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_Transconductor_26 out1 outVoltageBiasXXpXX2 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
m_FullyDifferential_SecondStage1_Transconductor_27 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_StageBias_28 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias nmos
m_FullyDifferential_SecondStage2_StageBias_29 SecondStage2YinnerStageBias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_Transconductor_30 out2 outVoltageBiasXXpXX2 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
m_FullyDifferential_SecondStage2_Transconductor_31 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_32 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_33 ibias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_34 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
m_FullyDifferential_SecondStage1_StageBias_35 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_36 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_12_11

