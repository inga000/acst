** Name: two_stage_single_output_op_amp_148_7

.MACRO two_stage_single_output_op_amp_148_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=30e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=258e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=297e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=42e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
mMainBias9 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=111e-6
mSecondStage1StageBias10 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=30e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=42e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=485e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=485e-6
mSimpleFirstStageLoad15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=526e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=382e-6
mSimpleFirstStageLoad17 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=526e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.5e-12
.EOM two_stage_single_output_op_amp_148_7

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 6.74601 mW
** Area: 5938 (mu_m)^2
** Transit frequency: 5.66901 MHz
** Transit frequency with error factor: 5.66547 MHz
** Slew rate: 6.79443 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** VoutMax: 4.67001 V
** VoutMin: 0.210001 V
** VcmMax: 5.09001 V
** VcmMin: 0.810001 V


** Expected Currents: 
** NormalTransistorNmos: 1.38963e+08 muA
** DiodeTransistorNmos: 1.79919e+08 muA
** DiodeTransistorNmos: 1.79918e+08 muA
** NormalTransistorNmos: 1.79917e+08 muA
** NormalTransistorNmos: 1.79918e+08 muA
** NormalTransistorPmos: -2.23039e+08 muA
** NormalTransistorPmos: -2.23038e+08 muA
** NormalTransistorPmos: -2.23037e+08 muA
** NormalTransistorPmos: -2.23038e+08 muA
** NormalTransistorNmos: 8.62431e+07 muA
** NormalTransistorNmos: 4.31211e+07 muA
** NormalTransistorNmos: 4.31211e+07 muA
** NormalTransistorNmos: 7.54155e+08 muA
** NormalTransistorPmos: -7.54154e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.38962e+08 muA
** DiodeTransistorPmos: -1.38961e+08 muA


** Expected Voltages: 
** ibias: 0.615001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.53801  V
** out: 2.5  V
** outFirstStage: 4.10201  V
** outSourceVoltageBiasXXpXX1: 4.27501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 1.15501  V
** innerTransistorStack1Load2: 4.25601  V
** innerTransistorStack2Load1: 1.15601  V
** innerTransistorStack2Load2: 4.25601  V
** out1: 2.09501  V
** sourceTransconductance: 1.90401  V


.END