** Name: two_stage_single_output_op_amp_64_8

.MACRO two_stage_single_output_op_amp_64_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=21e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=29e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=69e-6
mFoldedCascodeFirstStageLoad4 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=132e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=82e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=278e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerOutputLoad2 outInputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=27e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=27e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=254e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=130e-6
mFoldedCascodeFirstStageLoad12 outFirstStage outInputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=132e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=99e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=99e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=278e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=82e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=143e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=69e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=453e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.70001e-12
.EOM two_stage_single_output_op_amp_64_8

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 3.30901 mW
** Area: 10759 (mu_m)^2
** Transit frequency: 2.61401 MHz
** Transit frequency with error factor: 2.61418 MHz
** Slew rate: 5.08774 V/mu_s
** Phase margin: 60.1606°
** CMRR: 136 dB
** VoutMax: 4.25 V
** VoutMin: 0.760001 V
** VcmMax: 3.15001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -5.52349e+07 muA
** NormalTransistorNmos: 3.41991e+07 muA
** NormalTransistorNmos: 5.14251e+07 muA
** NormalTransistorNmos: 3.41991e+07 muA
** NormalTransistorNmos: 5.14251e+07 muA
** DiodeTransistorPmos: -3.41999e+07 muA
** DiodeTransistorPmos: -3.42009e+07 muA
** NormalTransistorPmos: -3.41999e+07 muA
** NormalTransistorPmos: -3.42009e+07 muA
** NormalTransistorPmos: -3.44549e+07 muA
** DiodeTransistorPmos: -3.44559e+07 muA
** NormalTransistorPmos: -1.72269e+07 muA
** NormalTransistorPmos: -1.72269e+07 muA
** NormalTransistorNmos: 4.83775e+08 muA
** NormalTransistorNmos: 4.83776e+08 muA
** NormalTransistorPmos: -4.83774e+08 muA
** DiodeTransistorNmos: 5.52341e+07 muA
** DiodeTransistorNmos: 5.52351e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.46401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.13601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.23301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 3.46501  V
** innerTransistorStack1Load2: 4.26501  V
** innerTransistorStack2Load2: 4.26401  V
** sourceGCC1: 0.529001  V
** sourceGCC2: 0.529001  V
** sourceTransconductance: 3.375  V
** innerStageBias: 0.521001  V
** inner: 4.23001  V


.END