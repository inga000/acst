.suckt  two_stage_fully_differential_op_amp_72_6 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outVoltageBiasXXpXX3 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_3 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_4 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_5 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_6 inputVoltageBiasXXnXX4 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_7 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_8 outFeedback outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX3 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m_FullyDifferential_FeedbackdStage_StageBias_10 FeedbackStageYinnerStageBias1 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_11 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX3 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m_FullyDifferential_FeedbackdStage_StageBias_12 FeedbackStageYinnerStageBias2 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackStage_Transconductor_13 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_14 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_15 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FeedbackStage_Transconductor_16 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FirstStage_Load_17 out1FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m_FullyDifferential_FirstStage_Load_18 out2FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m_FullyDifferential_FirstStage_Load_19 out1FirstStage outVoltageBiasXXpXX3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m_FullyDifferential_FirstStage_Load_20 FirstStageYinnerTransistorStack1Load2 outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_21 out2FirstStage outVoltageBiasXXpXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m_FullyDifferential_FirstStage_Load_22 FirstStageYinnerTransistorStack2Load2 outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_StageBias_23 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_FullyDifferential_FirstStage_StageBias_24 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Transconductor_25 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m_FullyDifferential_FirstStage_Transconductor_26 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_Transconductor_27 out1 inputVoltageBiasXXnXX3 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m_FullyDifferential_SecondStage1_Transconductor_28 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_29 out1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_FullyDifferential_SecondStage1_StageBias_30 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_Transconductor_31 out2 inputVoltageBiasXXnXX3 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m_FullyDifferential_SecondStage2_Transconductor_32 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_StageBias_33 out2 ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m_FullyDifferential_SecondStage2_StageBias_34 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_35 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_FullyDifferential_MainBias_36 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_37 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos
m_FullyDifferential_SecondStage1_StageBias_38 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_39 inputVoltageBiasXXnXX4 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_40 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_FullyDifferential_MainBias_41 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_42 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m_FullyDifferential_MainBias_43 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_44 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_72_6

