.suckt  complementary_op_amp9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 FirstStageYinnerOutputLoadNmos inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m4 FirstStageYinnerTransistorStack1LoadPmos outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m5 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m6 FirstStageYinnerTransistorStack2LoadPmos outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m7 FirstStageYinnerOutputLoadNmos FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m8 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos sourceNmos sourceNmos nmos
m9 out FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m10 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack1LoadNmos sourceNmos sourceNmos nmos
m11 FirstStageYsourceTransconductanceNmos ibias sourceNmos sourceNmos nmos
m12 FirstStageYsourceTransconductancePmos outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m13 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m14 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m15 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m16 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c1 out sourceNmos 
m17 ibias ibias sourceNmos sourceNmos nmos
m18 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m19 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end complementary_op_amp9

