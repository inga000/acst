** Name: two_stage_single_output_op_amp_57_12

.MACRO two_stage_single_output_op_amp_57_12 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=67e-6
m2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=14e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=290e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=12e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
m6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=19e-6
m7 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=55e-6
m8 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=290e-6
m9 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=24e-6
m10 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=9e-6
m11 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=24e-6
m12 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=17e-6
m13 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=17e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=67e-6
m15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=297e-6
m16 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=129e-6
m17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=541e-6
m18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=55e-6
m19 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=129e-6
m20 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=197e-6
m21 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=197e-6
m22 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=4e-6 W=596e-6
m23 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 7e-12
.EOM two_stage_single_output_op_amp_57_12

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 5.40901 mW
** Area: 14995 (mu_m)^2
** Transit frequency: 5.01801 MHz
** Transit frequency with error factor: 5.01119 MHz
** Slew rate: 8.30994 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** VoutMax: 4.25 V
** VoutMin: 1.12001 V
** VcmMax: 3.15001 V
** VcmMin: 0.0900001 V


** Expected Currents: 
** NormalTransistorNmos: 4.74531e+07 muA
** NormalTransistorPmos: -1.43135e+08 muA
** NormalTransistorPmos: -6.20209e+07 muA
** NormalTransistorNmos: 5.83331e+07 muA
** NormalTransistorNmos: 8.96341e+07 muA
** NormalTransistorNmos: 5.83331e+07 muA
** NormalTransistorNmos: 8.96341e+07 muA
** DiodeTransistorPmos: -5.83339e+07 muA
** NormalTransistorPmos: -5.83339e+07 muA
** NormalTransistorPmos: -6.26029e+07 muA
** NormalTransistorPmos: -6.26019e+07 muA
** NormalTransistorPmos: -3.13019e+07 muA
** NormalTransistorPmos: -3.13019e+07 muA
** NormalTransistorNmos: 6.30019e+08 muA
** DiodeTransistorNmos: 6.30018e+08 muA
** NormalTransistorPmos: -6.30018e+08 muA
** NormalTransistorPmos: -6.30019e+08 muA
** DiodeTransistorNmos: 1.43136e+08 muA
** NormalTransistorNmos: 1.43137e+08 muA
** DiodeTransistorNmos: 6.20201e+07 muA
** DiodeTransistorNmos: 6.20191e+07 muA
** DiodeTransistorPmos: -4.74539e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.15201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.52401  V
** inputVoltageBiasXXnXX2: 2.07001  V
** out: 2.5  V
** outFirstStage: 4.19401  V
** outSourceVoltageBiasXXnXX1: 0.762001  V
** outSourceVoltageBiasXXnXX2: 1.06201  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40301  V
** out1: 4.19201  V
** sourceGCC1: 1.21501  V
** sourceGCC2: 1.21501  V
** sourceTransconductance: 3.34601  V
** innerTransconductance: 4.75801  V
** inner: 0.763001  V


.END