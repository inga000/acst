** Name: two_stage_single_output_op_amp_100_2

.MACRO two_stage_single_output_op_amp_100_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=27e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=36e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
m5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=24e-6
m6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=127e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=591e-6
m8 inputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=342e-6
m9 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=193e-6
m10 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=36e-6
m11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=125e-6
m12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=194e-6
m13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=132e-6
m14 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=592e-6
m15 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=52e-6
m16 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
m17 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=591e-6
m18 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=52e-6
m19 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=63e-6
m20 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=63e-6
m21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=127e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_100_2

** Expected Performance Values: 
** Gain: 104 dB
** Power consumption: 3.45601 mW
** Area: 14243 (mu_m)^2
** Transit frequency: 9.77601 MHz
** Transit frequency with error factor: 9.7672 MHz
** Slew rate: 15.0209 V/mu_s
** Phase margin: 61.8795°
** CMRR: 96 dB
** VoutMax: 4.81001 V
** VoutMin: 0.300001 V
** VcmMax: 3 V
** VcmMin: 0.180001 V


** Expected Currents: 
** NormalTransistorNmos: 3.74031e+07 muA
** NormalTransistorNmos: 1.0359e+08 muA
** NormalTransistorPmos: -8.20499e+06 muA
** NormalTransistorPmos: -8.29749e+07 muA
** NormalTransistorPmos: -3.42849e+07 muA
** NormalTransistorPmos: -3.42849e+07 muA
** DiodeTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorPmos: -1.72162e+08 muA
** DiodeTransistorPmos: -1.72163e+08 muA
** NormalTransistorPmos: -3.42859e+07 muA
** NormalTransistorPmos: -3.42859e+07 muA
** NormalTransistorNmos: 3.70377e+08 muA
** NormalTransistorNmos: 3.70376e+08 muA
** NormalTransistorPmos: -3.70376e+08 muA
** DiodeTransistorNmos: 8.20401e+06 muA
** DiodeTransistorNmos: 8.29741e+07 muA
** DiodeTransistorPmos: -3.74039e+07 muA
** NormalTransistorPmos: -3.74049e+07 muA
** DiodeTransistorPmos: -1.03589e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXpXX2: 2.25701  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.24601  V
** outSourceVoltageBiasXXpXX1: 4.12201  V
** outVoltageBiasXXnXX0: 0.574001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.31001  V
** out1: 0.555001  V
** sourceGCC1: 3.01401  V
** sourceGCC2: 3.01301  V
** innerTransconductance: 0.150001  V
** inner: 4.12301  V


.END