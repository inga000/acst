** Name: two_stage_single_output_op_amp_6_4

.MACRO two_stage_single_output_op_amp_6_4 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=69e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=5e-6 W=69e-6
mSecondStage1StageBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias4 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=31e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=32e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=106e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=69e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=10e-6 W=214e-6
mSecondStage1Transconductor9 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=84e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=69e-6
mMainBias11 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=192e-6
mSimpleFirstStageTransconductor12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=23e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=170e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=529e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=561e-6
mSecondStage1StageBias16 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=413e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=23e-6
mMainBias18 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=548e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_6_4

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 8.33201 mW
** Area: 13376 (mu_m)^2
** Transit frequency: 2.79001 MHz
** Transit frequency with error factor: 2.77979 MHz
** Slew rate: 6.81262 V/mu_s
** Phase margin: 60.7336°
** CMRR: 93 dB
** negPSRR: 95 dB
** posPSRR: 132 dB
** VoutMax: 4.59001 V
** VoutMin: 0.460001 V
** VcmMax: 3.5 V
** VcmMin: 0.550001 V


** Expected Currents: 
** NormalTransistorNmos: 1.07627e+09 muA
** NormalTransistorPmos: -1.73659e+08 muA
** NormalTransistorPmos: -1.75041e+08 muA
** DiodeTransistorNmos: 2.69351e+07 muA
** NormalTransistorNmos: 2.69341e+07 muA
** NormalTransistorNmos: 2.69351e+07 muA
** DiodeTransistorNmos: 2.69341e+07 muA
** NormalTransistorPmos: -5.38719e+07 muA
** NormalTransistorPmos: -2.69359e+07 muA
** NormalTransistorPmos: -2.69359e+07 muA
** NormalTransistorNmos: 1.67638e+08 muA
** NormalTransistorNmos: 1.67637e+08 muA
** NormalTransistorPmos: -1.67637e+08 muA
** NormalTransistorPmos: -1.67638e+08 muA
** DiodeTransistorNmos: 1.7366e+08 muA
** DiodeTransistorNmos: 1.75042e+08 muA
** DiodeTransistorPmos: -1.07626e+09 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.862001  V
** out: 2.5  V
** outFirstStage: 0.709001  V
** outVoltageBiasXXnXX0: 1.08301  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.557001  V
** innerTransistorStack1Load1: 0.557001  V
** out1: 1.11401  V
** sourceTransconductance: 3.73801  V
** innerStageBias: 4.40001  V
** innerTransconductance: 0.304001  V


.END