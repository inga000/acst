** Name: two_stage_single_output_op_amp_138_3

.MACRO two_stage_single_output_op_amp_138_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=17e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=3e-6 W=9e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=9e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=9e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=127e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=127e-6
mSimpleFirstStageLoad9 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=112e-6
mMainBias10 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=14e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=160e-6
mSimpleFirstStageLoad12 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=112e-6
mMainBias13 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=35e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=3e-6 W=9e-6
mSimpleFirstStageTransconductor15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=50e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=61e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=479e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=500e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=9e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=50e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_138_3

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 2.03501 mW
** Area: 9424 (mu_m)^2
** Transit frequency: 3.26501 MHz
** Transit frequency with error factor: 3.25923 MHz
** Slew rate: 7.68636 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 0.350001 V
** VcmMax: 3.62001 V
** VcmMin: -0.25 V


** Expected Currents: 
** NormalTransistorNmos: 1.33331e+07 muA
** NormalTransistorNmos: 5.33601e+06 muA
** DiodeTransistorPmos: -3.04599e+07 muA
** NormalTransistorPmos: -3.04599e+07 muA
** NormalTransistorPmos: -3.04599e+07 muA
** DiodeTransistorPmos: -3.04599e+07 muA
** NormalTransistorNmos: 4.83771e+07 muA
** NormalTransistorNmos: 4.83781e+07 muA
** NormalTransistorNmos: 4.83771e+07 muA
** NormalTransistorNmos: 4.83781e+07 muA
** NormalTransistorPmos: -3.58369e+07 muA
** NormalTransistorPmos: -1.79179e+07 muA
** NormalTransistorPmos: -1.79179e+07 muA
** NormalTransistorNmos: 2.81665e+08 muA
** NormalTransistorPmos: -2.81664e+08 muA
** NormalTransistorPmos: -2.81665e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.33339e+07 muA
** DiodeTransistorPmos: -5.33699e+06 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.99201  V
** out: 2.5  V
** outFirstStage: 0.760001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.581001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.581001  V
** out1: 2.37201  V
** sourceTransconductance: 3.43701  V
** innerStageBias: 4.55601  V


.END