** Name: two_stage_single_output_op_amp_144_9

.MACRO two_stage_single_output_op_amp_144_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=4e-6 W=36e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=8e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=479e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=20e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=4e-6 W=36e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=479e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=71e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=20e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=435e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=435e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=599e-6
mMainBias17 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=393e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=599e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_144_9

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 7.99101 mW
** Area: 9402 (mu_m)^2
** Transit frequency: 3.62701 MHz
** Transit frequency with error factor: 3.62149 MHz
** Slew rate: 6.48337 V/mu_s
** Phase margin: 62.4525°
** CMRR: 120 dB
** VoutMax: 4.25 V
** VoutMin: 0.910001 V
** VcmMax: 4.97001 V
** VcmMin: 0.850001 V


** Expected Currents: 
** NormalTransistorPmos: -1.11209e+07 muA
** NormalTransistorPmos: -2.00229e+07 muA
** NormalTransistorNmos: 4.25806e+08 muA
** NormalTransistorNmos: 4.25807e+08 muA
** DiodeTransistorNmos: 4.25806e+08 muA
** NormalTransistorPmos: -4.41035e+08 muA
** NormalTransistorPmos: -4.41036e+08 muA
** NormalTransistorPmos: -4.41036e+08 muA
** NormalTransistorPmos: -4.41036e+08 muA
** NormalTransistorNmos: 3.04591e+07 muA
** NormalTransistorNmos: 1.52301e+07 muA
** NormalTransistorNmos: 1.52301e+07 muA
** NormalTransistorNmos: 6.65048e+08 muA
** DiodeTransistorNmos: 6.65047e+08 muA
** NormalTransistorPmos: -6.65047e+08 muA
** DiodeTransistorNmos: 1.11201e+07 muA
** NormalTransistorNmos: 1.11191e+07 muA
** DiodeTransistorNmos: 2.00221e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.32001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.660001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.562001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.17501  V
** innerTransistorStack2Load1: 1.15501  V
** innerTransistorStack2Load2: 4.17501  V
** out1: 2.09501  V
** sourceTransconductance: 1.81001  V
** inner: 0.658001  V


.END