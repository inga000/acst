** Name: one_stage_single_output_op_amp64

.MACRO one_stage_single_output_op_amp64 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=53e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=38e-6
m3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=68e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=511e-6
m5 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=10e-6
m6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=79e-6
m7 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=49e-6
m8 FirstStageYinnerOutputLoad2 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=49e-6
m9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
m10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
m11 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=390e-6
m12 out FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=10e-6
m13 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=79e-6
m14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=227e-6
m15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=227e-6
m16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=511e-6
m17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=68e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp64

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 1.46801 mW
** Area: 7171 (mu_m)^2
** Transit frequency: 3.60001 MHz
** Transit frequency with error factor: 3.60004 MHz
** Slew rate: 3.50003 V/mu_s
** Phase margin: 88.2356°
** CMRR: 129 dB
** VoutMax: 3.59001 V
** VoutMin: 0.860001 V
** VcmMax: 3.39001 V
** VcmMin: -0.329999 V


** Expected Currents: 
** NormalTransistorPmos: -5.76349e+07 muA
** NormalTransistorNmos: 7.00501e+07 muA
** NormalTransistorNmos: 1.07943e+08 muA
** NormalTransistorNmos: 7.00461e+07 muA
** NormalTransistorNmos: 1.07939e+08 muA
** DiodeTransistorPmos: -7.00489e+07 muA
** DiodeTransistorPmos: -7.00479e+07 muA
** NormalTransistorPmos: -7.00469e+07 muA
** NormalTransistorPmos: -7.00479e+07 muA
** NormalTransistorPmos: -7.57859e+07 muA
** DiodeTransistorPmos: -7.57849e+07 muA
** NormalTransistorPmos: -3.78929e+07 muA
** NormalTransistorPmos: -3.78929e+07 muA
** DiodeTransistorNmos: 5.76341e+07 muA
** DiodeTransistorNmos: 5.76351e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.55701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.23901  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.638001  V
** outSourceVoltageBiasXXpXX1: 4.27901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 3.02001  V
** innerTransistorStack1Load2: 4.21301  V
** innerTransistorStack2Load2: 4.20701  V
** sourceGCC1: 0.608001  V
** sourceGCC2: 0.608001  V
** sourceTransconductance: 3.23101  V
** inner: 4.27801  V


.END