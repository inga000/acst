** Name: two_stage_single_output_op_amp_196_12

.MACRO two_stage_single_output_op_amp_196_12 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=10e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=40e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=589e-6
m5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=149e-6
m6 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=8e-6 W=294e-6
m7 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
m8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=45e-6
m9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
m10 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=589e-6
m11 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=294e-6
m12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=30e-6
m13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=146e-6
m14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=149e-6
m15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=30e-6
m16 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=30e-6
m17 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=40e-6
m18 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
m19 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=500e-6
m20 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=286e-6
m21 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
m22 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=286e-6
m23 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=561e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 5.20001e-12
.EOM two_stage_single_output_op_amp_196_12

** Expected Performance Values: 
** Gain: 107 dB
** Power consumption: 12.8581 mW
** Area: 14991 (mu_m)^2
** Transit frequency: 5.67401 MHz
** Transit frequency with error factor: 5.52883 MHz
** Slew rate: 5.34706 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** VoutMax: 4.25 V
** VoutMin: 0.710001 V
** VcmMax: 4.81001 V
** VcmMin: 1.56001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00071e+07 muA
** NormalTransistorNmos: 1.43782e+08 muA
** NormalTransistorPmos: -3.83409e+07 muA
** DiodeTransistorNmos: 8.81599e+08 muA
** DiodeTransistorNmos: 8.81598e+08 muA
** NormalTransistorNmos: 8.81597e+08 muA
** NormalTransistorNmos: 8.81598e+08 muA
** NormalTransistorPmos: -8.95881e+08 muA
** NormalTransistorPmos: -8.95881e+08 muA
** NormalTransistorNmos: 2.85691e+07 muA
** DiodeTransistorNmos: 2.85681e+07 muA
** NormalTransistorNmos: 1.42851e+07 muA
** NormalTransistorNmos: 1.42851e+07 muA
** NormalTransistorNmos: 5.77795e+08 muA
** DiodeTransistorNmos: 5.77796e+08 muA
** NormalTransistorPmos: -5.77794e+08 muA
** NormalTransistorPmos: -5.77795e+08 muA
** DiodeTransistorNmos: 3.83401e+07 muA
** NormalTransistorNmos: 3.83391e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.00079e+07 muA
** DiodeTransistorPmos: -1.43781e+08 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.19501  V
** outInputVoltageBiasXXnXX1: 1.40901  V
** outSourceVoltageBiasXXnXX1: 0.705001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX2: 3.84101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack2Load1: 1.15601  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.75701  V
** inner: 0.702001  V
** inner: 0.556001  V


.END