** Name: two_stage_single_output_op_amp_195_8

.MACRO two_stage_single_output_op_amp_195_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=26e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
m3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=11e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=11e-6
m5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=9e-6
m6 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=301e-6
m7 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=11e-6
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=24e-6
m9 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=42e-6
m10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=120e-6
m11 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=11e-6
m12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=24e-6
m13 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=97e-6
m14 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
m15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=564e-6
m16 outFirstStage outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=59e-6
m17 FirstStageYout1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=59e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 13e-12
.EOM two_stage_single_output_op_amp_195_8

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 2.32101 mW
** Area: 7619 (mu_m)^2
** Transit frequency: 3.72401 MHz
** Transit frequency with error factor: 3.71298 MHz
** Slew rate: 3.5098 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** VoutMax: 4.85001 V
** VoutMin: 0.770001 V
** VcmMax: 4.70001 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorNmos: 1.61021e+07 muA
** DiodeTransistorNmos: 8.07651e+07 muA
** DiodeTransistorNmos: 8.07641e+07 muA
** NormalTransistorNmos: 8.07651e+07 muA
** NormalTransistorNmos: 8.07641e+07 muA
** NormalTransistorPmos: -1.03621e+08 muA
** NormalTransistorPmos: -1.03621e+08 muA
** NormalTransistorNmos: 4.57111e+07 muA
** NormalTransistorNmos: 4.57121e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.30865e+08 muA
** NormalTransistorNmos: 2.30864e+08 muA
** NormalTransistorPmos: -2.30864e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.61029e+07 muA


** Expected Voltages: 
** ibias: 1.11001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.28401  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 3.73201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.12901  V
** innerStageBias: 0.538001  V
** innerTransistorStack2Load1: 1.12901  V
** out1: 2.25901  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.492001  V


.END