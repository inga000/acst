.suckt  two_stage_single_output_op_amp_151_9 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
m5 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
m7 FirstStageYout1 ibias sourcePmos sourcePmos pmos
m8 outFirstStage ibias sourcePmos sourcePmos pmos
m9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c2 out sourceNmos 
m12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m13 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m14 out outFirstStage sourcePmos sourcePmos pmos
m15 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m16 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m17 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m18 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_151_9

