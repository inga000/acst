** Name: symmetrical_op_amp56

.MACRO symmetrical_op_amp56 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=28e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=28e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=21e-6
mSecondStage1StageBias5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=41e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=5e-6 W=41e-6
mSymmetricalFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=48e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=85e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=85e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=3e-6 W=19e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=19e-6
mSymmetricalFirstStageStageBias12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=48e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias13 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=41e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mMainBias15 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=95e-6
mSymmetricalFirstStageTransconductor16 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=16e-6
mSecondStage1StageBias17 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=5e-6 W=41e-6
mSymmetricalFirstStageTransconductor18 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=16e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp56

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 0.799001 mW
** Area: 3048 (mu_m)^2
** Transit frequency: 2.78601 MHz
** Transit frequency with error factor: 2.7862 MHz
** Slew rate: 3.5005 V/mu_s
** Phase margin: 68.755°
** CMRR: 143 dB
** negPSRR: 49 dB
** posPSRR: 57 dB
** VoutMax: 3.45001 V
** VoutMin: 0.430001 V
** VcmMax: 3.10001 V
** VcmMin: 0.0100001 V


** Expected Currents: 
** NormalTransistorPmos: -4.61019e+07 muA
** DiodeTransistorNmos: 1.16461e+07 muA
** DiodeTransistorNmos: 1.16461e+07 muA
** NormalTransistorPmos: -2.32949e+07 muA
** DiodeTransistorPmos: -2.32939e+07 muA
** NormalTransistorPmos: -1.16469e+07 muA
** NormalTransistorPmos: -1.16469e+07 muA
** NormalTransistorNmos: 3.50281e+07 muA
** NormalTransistorNmos: 3.50271e+07 muA
** NormalTransistorPmos: -3.50289e+07 muA
** DiodeTransistorPmos: -3.50299e+07 muA
** DiodeTransistorPmos: -3.54219e+07 muA
** NormalTransistorPmos: -3.54229e+07 muA
** NormalTransistorNmos: 3.54211e+07 muA
** NormalTransistorNmos: 3.54201e+07 muA
** DiodeTransistorNmos: 4.61011e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.30201  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.832001  V
** inSourceStageBiasComplementarySecondStage: 3.94501  V
** inSourceTransconductanceComplementarySecondStage: 0.576001  V
** innerComplementarySecondStage: 2.89001  V
** out: 2.5  V
** outFirstStage: 0.576001  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.26501  V
** innerTransconductance: 0.171001  V
** inner: 3.94401  V
** inner: 0.171001  V
** inner: 4.14801  V


.END