** Name: symmetrical_op_amp9

.MACRO symmetrical_op_amp9 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=19e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSymmetricalFirstStageLoad4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=19e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=61e-6
mMainBias6 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
mMainBias9 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=3e-6 W=36e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=36e-6
mSymmetricalFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=5e-6 W=439e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=42e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias14 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=42e-6
mMainBias15 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=5e-6 W=89e-6
mSymmetricalFirstStageTransconductor16 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=166e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias17 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=3e-6 W=75e-6
mMainBias18 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=15e-6
mSecondStage1StageBias19 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=335e-6
mSymmetricalFirstStageTransconductor20 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=166e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp9

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 1.07501 mW
** Area: 6256 (mu_m)^2
** Transit frequency: 3.28001 MHz
** Transit frequency with error factor: 3.28048 MHz
** Slew rate: 4.55319 V/mu_s
** Phase margin: 88.2356°
** CMRR: 150 dB
** negPSRR: 49 dB
** posPSRR: 58 dB
** VoutMax: 4.42001 V
** VoutMin: 0.360001 V
** VcmMax: 4 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 1.32801e+07 muA
** NormalTransistorPmos: -2.50299e+06 muA
** NormalTransistorPmos: -1.48519e+07 muA
** DiodeTransistorNmos: 3.61881e+07 muA
** DiodeTransistorNmos: 3.61881e+07 muA
** NormalTransistorPmos: -7.23789e+07 muA
** NormalTransistorPmos: -3.61889e+07 muA
** NormalTransistorPmos: -3.61889e+07 muA
** NormalTransistorNmos: 4.57111e+07 muA
** NormalTransistorNmos: 4.57121e+07 muA
** NormalTransistorPmos: -4.57119e+07 muA
** NormalTransistorPmos: -4.57129e+07 muA
** NormalTransistorPmos: -4.61739e+07 muA
** NormalTransistorPmos: -4.61749e+07 muA
** NormalTransistorNmos: 4.61731e+07 muA
** NormalTransistorNmos: 4.61721e+07 muA
** DiodeTransistorNmos: 2.50201e+06 muA
** DiodeTransistorNmos: 1.48511e+07 muA
** DiodeTransistorPmos: -1.32809e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.22101  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 3.68601  V
** inOutputTransconductanceComplementarySecondStage: 0.768001  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 4.00701  V
** inputVoltageBiasXXnXX0: 0.577001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.28401  V
** innerStageBias: 4.40101  V
** innerTransconductance: 0.150001  V
** inner: 4.57001  V
** inner: 0.150001  V


.END