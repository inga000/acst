.suckt  one_stage_single_output_op_amp9 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m2 out FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos
m3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m6 out in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m7 ibias ibias sourceNmos sourceNmos nmos
.end one_stage_single_output_op_amp9

