** Name: two_stage_single_output_op_amp_29_7

.MACRO two_stage_single_output_op_amp_29_7 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
m3 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=21e-6
m4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
m5 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
m6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=18e-6
m7 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m8 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=41e-6
m9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=18e-6
m10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=91e-6
m11 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=48e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=293e-6
m13 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_29_7

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 5.55801 mW
** Area: 3156 (mu_m)^2
** Transit frequency: 7.98201 MHz
** Transit frequency with error factor: 7.9719 MHz
** Slew rate: 7.52287 V/mu_s
** Phase margin: 60.1606°
** CMRR: 94 dB
** negPSRR: 158 dB
** posPSRR: 92 dB
** VoutMax: 4.56001 V
** VoutMin: 0.200001 V
** VcmMax: 4.40001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorNmos: 8.21501e+06 muA
** NormalTransistorPmos: -1.91489e+07 muA
** DiodeTransistorPmos: -3.42849e+07 muA
** NormalTransistorPmos: -3.42849e+07 muA
** NormalTransistorNmos: 6.85671e+07 muA
** NormalTransistorNmos: 6.85661e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 1.00565e+09 muA
** NormalTransistorPmos: -1.00564e+09 muA
** DiodeTransistorNmos: 1.91481e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.21599e+06 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.879001  V
** out: 2.5  V
** outFirstStage: 3.99601  V
** outVoltageBiasXXpXX0: 3.99001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.242001  V
** out1: 3.99601  V
** sourceTransconductance: 1.94501  V


.END