.suckt  symmetrical_op_amp71 ibias in1 in2 out sourceNmos sourcePmos
m1 outFirstStage outFirstStage sourcePmos sourcePmos pmos
m2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m3 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m5 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m6 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m7 out innerComplementarySecondStage sourceNmos sourceNmos nmos
m8 out outFirstStage sourcePmos sourcePmos pmos
m9 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
m10 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m11 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
.end symmetrical_op_amp71

