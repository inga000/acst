** Name: two_stage_single_output_op_amp_71_2

.MACRO two_stage_single_output_op_amp_71_2 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=22e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=256e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
m5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=68e-6
m6 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=110e-6
m7 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=477e-6
m8 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=256e-6
m9 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=43e-6
m10 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=52e-6
m11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=113e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=113e-6
m13 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=90e-6
m14 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=239e-6
m15 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=314e-6
m16 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=444e-6
m17 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=37e-6
m18 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=37e-6
m19 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=100e-6
m20 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=100e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 11.2001e-12
.EOM two_stage_single_output_op_amp_71_2

** Expected Performance Values: 
** Gain: 105 dB
** Power consumption: 6.29901 mW
** Area: 8906 (mu_m)^2
** Transit frequency: 8.08301 MHz
** Transit frequency with error factor: 8.07807 MHz
** Slew rate: 5.35473 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** VoutMax: 4.76001 V
** VoutMin: 0.300001 V
** VcmMax: 5.16001 V
** VcmMin: 1.35001 V


** Expected Currents: 
** NormalTransistorNmos: 1.82761e+08 muA
** NormalTransistorNmos: 7.12891e+07 muA
** NormalTransistorPmos: -3.23104e+08 muA
** NormalTransistorPmos: -6.05089e+07 muA
** NormalTransistorPmos: -1.03554e+08 muA
** NormalTransistorPmos: -6.05089e+07 muA
** NormalTransistorPmos: -1.03554e+08 muA
** DiodeTransistorNmos: 6.05081e+07 muA
** NormalTransistorNmos: 6.05081e+07 muA
** NormalTransistorNmos: 8.60891e+07 muA
** NormalTransistorNmos: 8.60881e+07 muA
** NormalTransistorNmos: 4.30451e+07 muA
** NormalTransistorNmos: 4.30451e+07 muA
** NormalTransistorNmos: 4.65485e+08 muA
** NormalTransistorNmos: 4.65484e+08 muA
** NormalTransistorPmos: -4.65484e+08 muA
** DiodeTransistorNmos: 3.23105e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.8276e+08 muA
** DiodeTransistorPmos: -7.12899e+07 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.997001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.556001  V
** outVoltageBiasXXpXX2: 4.19501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.442001  V
** out1: 0.563001  V
** sourceGCC1: 4.55101  V
** sourceGCC2: 4.55101  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 0.440001  V


.END