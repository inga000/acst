** Name: two_stage_single_output_op_amp_113_8

.MACRO two_stage_single_output_op_amp_113_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=7e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=12e-6
m3 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
m4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=59e-6
m6 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=211e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=18e-6
m8 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=25e-6
m9 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=57e-6
m10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=161e-6
m11 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=18e-6
m12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=127e-6
m13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=127e-6
m14 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
m15 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=33e-6
m16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=536e-6
m17 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=59e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_113_8

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 3.97601 mW
** Area: 4824 (mu_m)^2
** Transit frequency: 8.04001 MHz
** Transit frequency with error factor: 8.03505 MHz
** Slew rate: 17.503 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.75 V
** VoutMin: 0.820001 V
** VcmMax: 4.43001 V
** VcmMin: 1.37001 V


** Expected Currents: 
** NormalTransistorNmos: 2.50191e+07 muA
** NormalTransistorPmos: -9.05179e+07 muA
** NormalTransistorNmos: 3.45551e+07 muA
** NormalTransistorNmos: 3.45551e+07 muA
** DiodeTransistorPmos: -3.45559e+07 muA
** NormalTransistorPmos: -3.45559e+07 muA
** NormalTransistorNmos: 1.59629e+08 muA
** NormalTransistorNmos: 1.59628e+08 muA
** NormalTransistorNmos: 3.45561e+07 muA
** NormalTransistorNmos: 3.45561e+07 muA
** NormalTransistorNmos: 6.00478e+08 muA
** NormalTransistorNmos: 6.00477e+08 muA
** NormalTransistorPmos: -6.00477e+08 muA
** DiodeTransistorNmos: 9.05171e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.50199e+07 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.65001  V
** out: 2.5  V
** outFirstStage: 4.18501  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXpXX0: 3.88001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.483001  V
** out1: 4.17901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.481001  V


.END