** Name: one_stage_single_output_op_amp68

.MACRO one_stage_single_output_op_amp68 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=30e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=37e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=11e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=67e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=465e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=48e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=48e-6
mFoldedCascodeFirstStageLoad10 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=74e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=74e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=465e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=67e-6
mMainBias16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=534e-6
mFoldedCascodeFirstStageLoad17 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=11e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp68

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 1.54701 mW
** Area: 6787 (mu_m)^2
** Transit frequency: 3.42301 MHz
** Transit frequency with error factor: 3.42341 MHz
** Slew rate: 3.50001 V/mu_s
** Phase margin: 89.9544°
** CMRR: 130 dB
** VoutMax: 3.24001 V
** VoutMin: 0.770001 V
** VcmMax: 3.34001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorPmos: -7.93869e+07 muA
** NormalTransistorNmos: 7.00261e+07 muA
** NormalTransistorNmos: 1.0504e+08 muA
** NormalTransistorNmos: 7.00221e+07 muA
** NormalTransistorNmos: 1.05036e+08 muA
** DiodeTransistorPmos: -7.00249e+07 muA
** NormalTransistorPmos: -7.00239e+07 muA
** NormalTransistorPmos: -7.00229e+07 muA
** DiodeTransistorPmos: -7.00239e+07 muA
** NormalTransistorPmos: -7.00289e+07 muA
** DiodeTransistorPmos: -7.00299e+07 muA
** NormalTransistorPmos: -3.50139e+07 muA
** NormalTransistorPmos: -3.50139e+07 muA
** DiodeTransistorNmos: 7.93861e+07 muA
** DiodeTransistorNmos: 7.93871e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.50501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.14601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.565001  V
** outSourceVoltageBiasXXpXX1: 4.25301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 3.83201  V
** innerTransistorStack2Load2: 3.83701  V
** out1: 2.67401  V
** sourceGCC1: 0.537001  V
** sourceGCC2: 0.537001  V
** sourceTransconductance: 3.22601  V
** inner: 4.25101  V


.END