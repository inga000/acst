** Name: two_stage_single_output_op_amp_58_2

.MACRO two_stage_single_output_op_amp_58_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=80e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=65e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=582e-6
m6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=253e-6
m7 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=600e-6
m8 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=568e-6
m9 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=32e-6
m10 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=568e-6
m11 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=426e-6
m12 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=426e-6
m13 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=520e-6
m14 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=91e-6
m15 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=587e-6
m16 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=253e-6
m17 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=32e-6
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=130e-6
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=130e-6
m20 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=582e-6
m21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 14.9001e-12
.EOM two_stage_single_output_op_amp_58_2

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 7.30801 mW
** Area: 14982 (mu_m)^2
** Transit frequency: 5.25801 MHz
** Transit frequency with error factor: 5.24313 MHz
** Slew rate: 14.1123 V/mu_s
** Phase margin: 60.1606°
** CMRR: 88 dB
** VoutMax: 4.69001 V
** VoutMin: 0.350001 V
** VcmMax: 3.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorPmos: -2.67209e+07 muA
** NormalTransistorPmos: -7.61869e+07 muA
** NormalTransistorNmos: 2.70458e+08 muA
** NormalTransistorNmos: 4.06026e+08 muA
** NormalTransistorNmos: 2.70458e+08 muA
** NormalTransistorNmos: 4.06026e+08 muA
** DiodeTransistorPmos: -2.70457e+08 muA
** NormalTransistorPmos: -2.70457e+08 muA
** NormalTransistorPmos: -2.71138e+08 muA
** DiodeTransistorPmos: -2.71139e+08 muA
** NormalTransistorPmos: -1.35568e+08 muA
** NormalTransistorPmos: -1.35568e+08 muA
** NormalTransistorNmos: 4.96068e+08 muA
** NormalTransistorNmos: 4.96067e+08 muA
** NormalTransistorPmos: -4.96065e+08 muA
** DiodeTransistorNmos: 2.67201e+07 muA
** DiodeTransistorNmos: 7.61861e+07 muA
** DiodeTransistorPmos: -3.04759e+07 muA
** NormalTransistorPmos: -3.04769e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.54801  V
** outSourceVoltageBiasXXpXX1: 4.27401  V
** outVoltageBiasXXnXX1: 0.905001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.08901  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.60201  V
** innerTransconductance: 0.302001  V
** inner: 4.27401  V


.END