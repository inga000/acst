** Name: two_stage_single_output_op_amp_170_5

.MACRO two_stage_single_output_op_amp_170_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=22e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=6e-6 W=21e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=6e-6 W=21e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=13e-6
mMainBias6 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=139e-6
mSecondStage1StageBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=268e-6
mSimpleFirstStageLoad9 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=197e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=219e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=219e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=134e-6
mSimpleFirstStageLoad13 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=197e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
mMainBias15 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=139e-6
mSimpleFirstStageTransconductor16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=161e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=6e-6 W=21e-6
mSimpleFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=139e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mMainBias20 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=268e-6
mSimpleFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=6e-6 W=21e-6
mSimpleFirstStageTransconductor23 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=161e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.40001e-12
.EOM two_stage_single_output_op_amp_170_5

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 7.12301 mW
** Area: 10982 (mu_m)^2
** Transit frequency: 4.84001 MHz
** Transit frequency with error factor: 4.83687 MHz
** Slew rate: 10.4865 V/mu_s
** Phase margin: 60.1606°
** CMRR: 85 dB
** VoutMax: 3.43001 V
** VoutMin: 0.330001 V
** VcmMax: 3.20001 V
** VcmMin: -0.25 V


** Expected Currents: 
** NormalTransistorNmos: 6.37001e+06 muA
** NormalTransistorNmos: 4.47641e+07 muA
** DiodeTransistorPmos: -3.55359e+07 muA
** DiodeTransistorPmos: -3.55359e+07 muA
** NormalTransistorPmos: -3.55359e+07 muA
** NormalTransistorPmos: -3.55359e+07 muA
** NormalTransistorNmos: 6.97511e+07 muA
** NormalTransistorNmos: 6.97521e+07 muA
** NormalTransistorNmos: 6.97511e+07 muA
** NormalTransistorNmos: 6.97521e+07 muA
** NormalTransistorPmos: -6.84329e+07 muA
** DiodeTransistorPmos: -6.84339e+07 muA
** NormalTransistorPmos: -3.42159e+07 muA
** NormalTransistorPmos: -3.42159e+07 muA
** NormalTransistorNmos: 1.22394e+09 muA
** NormalTransistorPmos: -1.22393e+09 muA
** DiodeTransistorPmos: -1.22393e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -6.37099e+06 muA
** NormalTransistorPmos: -6.37199e+06 muA
** DiodeTransistorPmos: -4.47649e+07 muA
** NormalTransistorPmos: -4.47659e+07 muA


** Expected Voltages: 
** ibias: 1.14001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.735001  V
** outInputVoltageBiasXXpXX1: 3.54001  V
** outInputVoltageBiasXXpXX2: 2.86101  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outSourceVoltageBiasXXpXX1: 4.27001  V
** outSourceVoltageBiasXXpXX2: 3.93301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.576001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.576001  V
** sourceTransconductance: 3.40801  V
** inner: 4.26901  V
** inner: 3.92301  V


.END