.suckt  symmetrical_op_amp19 ibias in1 in2 out sourceNmos sourcePmos
m1 outFirstStage outFirstStage sourcePmos sourcePmos pmos
m2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m3 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m4 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m5 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m6 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m7 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
m8 out outFirstStage sourcePmos sourcePmos pmos
m9 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos
m10 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos
m11 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m12 ibias ibias sourceNmos sourceNmos nmos
.end symmetrical_op_amp19

