** Name: one_stage_single_output_op_amp59

.MACRO one_stage_single_output_op_amp59 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=18e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=35e-6
m3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=174e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=16e-6
m5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=10e-6 W=177e-6
m6 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=35e-6
m7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=35e-6
m8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=136e-6
m9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=136e-6
m10 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=3e-6 W=34e-6
m11 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=42e-6
m12 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=110e-6
m13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=10e-6 W=177e-6
m14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=346e-6
m15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=346e-6
m16 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=7e-6 W=599e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp59

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 1.28401 mW
** Area: 14972 (mu_m)^2
** Transit frequency: 3.70101 MHz
** Transit frequency with error factor: 3.70063 MHz
** Slew rate: 3.5004 V/mu_s
** Phase margin: 87.0896°
** CMRR: 128 dB
** VoutMax: 3.37001 V
** VoutMin: 0.960001 V
** VcmMax: 3.01001 V
** VcmMin: -0.349999 V


** Expected Currents: 
** NormalTransistorPmos: -2.66179e+07 muA
** NormalTransistorNmos: 7.00671e+07 muA
** NormalTransistorNmos: 1.051e+08 muA
** NormalTransistorNmos: 7.00681e+07 muA
** NormalTransistorNmos: 1.05101e+08 muA
** NormalTransistorPmos: -7.00679e+07 muA
** NormalTransistorPmos: -7.00689e+07 muA
** DiodeTransistorPmos: -7.00679e+07 muA
** NormalTransistorPmos: -7.00649e+07 muA
** NormalTransistorPmos: -7.00639e+07 muA
** NormalTransistorPmos: -3.50329e+07 muA
** NormalTransistorPmos: -3.50329e+07 muA
** DiodeTransistorNmos: 2.66171e+07 muA
** DiodeTransistorNmos: 2.66181e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.22501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.31801  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.618001  V
** outSourceVoltageBiasXXpXX1: 3.93901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 3.96301  V
** innerStageBias: 4.00201  V
** out1: 2.80801  V
** sourceGCC1: 0.568001  V
** sourceGCC2: 0.568001  V
** sourceTransconductance: 3.21401  V


.END