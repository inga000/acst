** Name: two_stage_single_output_op_amp_60_8

.MACRO two_stage_single_output_op_amp_60_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=12e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=8e-6 W=158e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=527e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=21e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=21e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=248e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=133e-6
mFoldedCascodeFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=28e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=28e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=8e-6 W=527e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=158e-6
mMainBias17 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=393e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=97e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=18e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.20001e-12
.EOM two_stage_single_output_op_amp_60_8

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 3.04501 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 2.72901 MHz
** Transit frequency with error factor: 2.729 MHz
** Slew rate: 3.82987 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 4.25 V
** VoutMin: 0.760001 V
** VcmMax: 3.22001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.48429e+07 muA
** NormalTransistorNmos: 2.37731e+07 muA
** NormalTransistorNmos: 4.07551e+07 muA
** NormalTransistorNmos: 2.37701e+07 muA
** NormalTransistorNmos: 4.07501e+07 muA
** NormalTransistorPmos: -2.37719e+07 muA
** NormalTransistorPmos: -2.37709e+07 muA
** DiodeTransistorPmos: -2.37719e+07 muA
** NormalTransistorPmos: -3.39619e+07 muA
** DiodeTransistorPmos: -3.39609e+07 muA
** NormalTransistorPmos: -1.69809e+07 muA
** NormalTransistorPmos: -1.69809e+07 muA
** NormalTransistorNmos: 4.8269e+08 muA
** NormalTransistorNmos: 4.82689e+08 muA
** NormalTransistorPmos: -4.82689e+08 muA
** DiodeTransistorNmos: 2.48421e+07 muA
** DiodeTransistorNmos: 2.48431e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.53301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11701  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outSourceVoltageBiasXXpXX1: 4.26701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.20001  V
** out1: 3.36301  V
** sourceGCC1: 0.544001  V
** sourceGCC2: 0.544001  V
** sourceTransconductance: 3.38201  V
** innerStageBias: 0.504001  V
** inner: 4.26501  V


.END