** Name: two_stage_single_output_op_amp_40_8

.MACRO two_stage_single_output_op_amp_40_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=8e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=377e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=181e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
m5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=139e-6
m6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=72e-6
m7 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=72e-6
m8 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=77e-6
m9 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=242e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=61e-6
m11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=61e-6
m12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=181e-6
m13 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=377e-6
m15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=350e-6
m16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=72e-6
m17 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=220e-6
m18 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=72e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_40_8

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 4.32501 mW
** Area: 13364 (mu_m)^2
** Transit frequency: 6.74501 MHz
** Transit frequency with error factor: 6.74102 MHz
** Slew rate: 6.35687 V/mu_s
** Phase margin: 60.1606°
** CMRR: 110 dB
** negPSRR: 109 dB
** posPSRR: 102 dB
** VoutMax: 4.69001 V
** VoutMin: 0.800001 V
** VcmMax: 3.98001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 7.68371e+07 muA
** NormalTransistorPmos: -1.1958e+08 muA
** DiodeTransistorPmos: -2.90469e+07 muA
** NormalTransistorPmos: -2.90479e+07 muA
** NormalTransistorPmos: -2.90469e+07 muA
** DiodeTransistorPmos: -2.90479e+07 muA
** NormalTransistorNmos: 5.80911e+07 muA
** DiodeTransistorNmos: 5.80901e+07 muA
** NormalTransistorNmos: 2.90461e+07 muA
** NormalTransistorNmos: 2.90461e+07 muA
** NormalTransistorNmos: 6.00478e+08 muA
** NormalTransistorNmos: 6.00477e+08 muA
** NormalTransistorPmos: -6.00477e+08 muA
** DiodeTransistorNmos: 1.19581e+08 muA
** NormalTransistorNmos: 1.19581e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.68379e+07 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.08601  V
** out: 2.5  V
** outFirstStage: 4.125  V
** outInputVoltageBiasXXnXX1: 1.15801  V
** outSourceVoltageBiasXXnXX1: 0.579001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.28501  V
** innerTransistorStack1Load1: 4.28401  V
** out1: 3.57001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.486001  V
** inner: 0.579001  V


.END