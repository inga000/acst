** Name: two_stage_single_output_op_amp_53_5

.MACRO two_stage_single_output_op_amp_53_5 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=31e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=3e-6 W=87e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=27e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=18e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=63e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=251e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=354e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=31e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=24e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=24e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=157e-6
mMainBias12 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=495e-6
mSecondStage1Transconductor13 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=169e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=87e-6
mMainBias15 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=506e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=92e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=164e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=164e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=63e-6
mSecondStage1StageBias20 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=251e-6
mFoldedCascodeFirstStageLoad21 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=92e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5e-12
.EOM two_stage_single_output_op_amp_53_5

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 6.38601 mW
** Area: 12082 (mu_m)^2
** Transit frequency: 5.38601 MHz
** Transit frequency with error factor: 5.38574 MHz
** Slew rate: 10.9315 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 3.63001 V
** VoutMin: 0.600001 V
** VcmMax: 5.24001 V
** VcmMin: 0.920001 V


** Expected Currents: 
** NormalTransistorNmos: 1.8554e+08 muA
** NormalTransistorNmos: 1.82761e+08 muA
** NormalTransistorPmos: -5.52359e+07 muA
** NormalTransistorPmos: -8.40209e+07 muA
** NormalTransistorPmos: -5.52359e+07 muA
** NormalTransistorPmos: -8.40209e+07 muA
** DiodeTransistorNmos: 5.52351e+07 muA
** DiodeTransistorNmos: 5.52341e+07 muA
** NormalTransistorNmos: 5.52351e+07 muA
** NormalTransistorNmos: 5.52341e+07 muA
** NormalTransistorNmos: 5.75691e+07 muA
** NormalTransistorNmos: 2.87841e+07 muA
** NormalTransistorNmos: 2.87841e+07 muA
** NormalTransistorNmos: 7.30877e+08 muA
** NormalTransistorPmos: -7.30876e+08 muA
** DiodeTransistorPmos: -7.30877e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.85539e+08 muA
** NormalTransistorPmos: -1.8554e+08 muA
** DiodeTransistorPmos: -1.8276e+08 muA
** DiodeTransistorPmos: -1.82761e+08 muA


** Expected Voltages: 
** ibias: 0.580001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.95201  V
** out: 2.5  V
** outFirstStage: 1.00601  V
** outInputVoltageBiasXXpXX1: 3.06201  V
** outSourceVoltageBiasXXpXX1: 4.03101  V
** outSourceVoltageBiasXXpXX2: 4.26601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.656001  V
** innerTransistorStack2Load2: 0.656001  V
** out1: 1.21101  V
** sourceGCC1: 3.69901  V
** sourceGCC2: 3.69901  V
** sourceTransconductance: 1.75701  V
** inner: 4.03001  V


.END