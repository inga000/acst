** Name: two_stage_single_output_op_amp_190_8

.MACRO two_stage_single_output_op_amp_190_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=45e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=28e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=22e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=138e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=42e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=9e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=10e-6
mSimpleFirstStageLoad9 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=45e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=138e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=173e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=28e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=180e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=10e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=243e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=243e-6
mSimpleFirstStageLoad18 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=600e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=119e-6
mSimpleFirstStageLoad20 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=600e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=13e-6
mMainBias22 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_190_8

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 6.15501 mW
** Area: 10433 (mu_m)^2
** Transit frequency: 3.75201 MHz
** Transit frequency with error factor: 3.74065 MHz
** Slew rate: 14.4505 V/mu_s
** Phase margin: 60.1606°
** CMRR: 102 dB
** VoutMax: 4.25 V
** VoutMin: 0.810001 V
** VcmMax: 4.59001 V
** VcmMin: 1.77001 V


** Expected Currents: 
** NormalTransistorPmos: -1.44989e+07 muA
** NormalTransistorPmos: -4.19029e+07 muA
** NormalTransistorNmos: 2.39891e+08 muA
** NormalTransistorNmos: 2.39892e+08 muA
** DiodeTransistorNmos: 2.39891e+08 muA
** NormalTransistorPmos: -2.75239e+08 muA
** NormalTransistorPmos: -2.75238e+08 muA
** NormalTransistorPmos: -2.75239e+08 muA
** NormalTransistorPmos: -2.75238e+08 muA
** NormalTransistorNmos: 7.06971e+07 muA
** DiodeTransistorNmos: 7.06961e+07 muA
** NormalTransistorNmos: 3.53491e+07 muA
** NormalTransistorNmos: 3.53491e+07 muA
** NormalTransistorNmos: 6.04127e+08 muA
** NormalTransistorNmos: 6.04126e+08 muA
** NormalTransistorPmos: -6.04126e+08 muA
** DiodeTransistorNmos: 1.44981e+07 muA
** NormalTransistorNmos: 1.44971e+07 muA
** DiodeTransistorNmos: 4.19021e+07 muA
** DiodeTransistorNmos: 4.19011e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.14001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.15801  V
** outInputVoltageBiasXXnXX2: 1.16301  V
** outSourceVoltageBiasXXnXX1: 0.579001  V
** outSourceVoltageBiasXXnXX2: 0.608001  V
** outSourceVoltageBiasXXpXX1: 3.93501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.02301  V
** innerTransistorStack2Load1: 1.15501  V
** innerTransistorStack2Load2: 4.02301  V
** out1: 2.09501  V
** sourceTransconductance: 1.47901  V
** innerStageBias: 0.558001  V
** inner: 0.578001  V


.END