** Name: two_stage_single_output_op_amp_104_7

.MACRO two_stage_single_output_op_amp_104_7 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=57e-6
m2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=152e-6
m4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=40e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=484e-6
m6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=10e-6
m7 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
m8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=174e-6
m9 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
m10 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=152e-6
m11 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=215e-6
m12 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=320e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=191e-6
m14 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=103e-6
m15 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=484e-6
m16 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=103e-6
m17 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=135e-6
m18 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=135e-6
m19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10.4001e-12
.EOM two_stage_single_output_op_amp_104_7

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 11.2391 mW
** Area: 13545 (mu_m)^2
** Transit frequency: 3.93701 MHz
** Transit frequency with error factor: 3.93689 MHz
** Slew rate: 11.716 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 3.47001 V
** VoutMin: 0.200001 V
** VcmMax: 3.08001 V
** VcmMin: 0.290001 V


** Expected Currents: 
** NormalTransistorNmos: 3.92501e+07 muA
** NormalTransistorPmos: -5.37459e+07 muA
** NormalTransistorPmos: -8.04939e+07 muA
** NormalTransistorPmos: -4.17159e+07 muA
** NormalTransistorPmos: -4.17149e+07 muA
** DiodeTransistorNmos: 4.17151e+07 muA
** NormalTransistorNmos: 4.17141e+07 muA
** NormalTransistorNmos: 4.17151e+07 muA
** NormalTransistorPmos: -1.22679e+08 muA
** DiodeTransistorPmos: -1.22678e+08 muA
** NormalTransistorPmos: -4.17149e+07 muA
** NormalTransistorPmos: -4.17149e+07 muA
** NormalTransistorNmos: 1.97086e+09 muA
** NormalTransistorPmos: -1.97085e+09 muA
** DiodeTransistorNmos: 5.37451e+07 muA
** DiodeTransistorNmos: 8.04931e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -3.92509e+07 muA


** Expected Voltages: 
** ibias: 3.39601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXnXX2: 0.601001  V
** out: 2.5  V
** outFirstStage: 2.90901  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXpXX2: 2.35001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.38501  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.06401  V
** sourceGCC2: 3.06401  V
** inner: 4.19601  V


.END