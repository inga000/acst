** Name: one_stage_single_output_op_amp87

.MACRO one_stage_single_output_op_amp87 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=140e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=29e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=24e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=4e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=140e-6
mTelescopicFirstStageLoad7 out inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=93e-6
mMainBias8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=12e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=357e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=206e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=206e-6
mMainBias12 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=55e-6
mTelescopicFirstStageLoad13 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=357e-6
mMainBias14 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=431e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp87

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 1.16801 mW
** Area: 6281 (mu_m)^2
** Transit frequency: 9.07001 MHz
** Transit frequency with error factor: 9.0699 MHz
** Slew rate: 9.04866 V/mu_s
** Phase margin: 64.7443°
** CMRR: 152 dB
** VoutMax: 4.34001 V
** VoutMin: 0.300001 V
** VcmMax: 4.02001 V
** VcmMin: 0.380001 V


** Expected Currents: 
** NormalTransistorNmos: 3.44301e+06 muA
** NormalTransistorPmos: -8.43799e+06 muA
** NormalTransistorPmos: -2.30869e+07 muA
** NormalTransistorPmos: -8.93339e+07 muA
** NormalTransistorPmos: -8.93349e+07 muA
** DiodeTransistorNmos: 8.93331e+07 muA
** NormalTransistorNmos: 8.93341e+07 muA
** NormalTransistorNmos: 8.93331e+07 muA
** NormalTransistorPmos: -1.8211e+08 muA
** NormalTransistorPmos: -8.93339e+07 muA
** NormalTransistorPmos: -8.93339e+07 muA
** DiodeTransistorNmos: 8.43701e+06 muA
** DiodeTransistorNmos: 2.30861e+07 muA
** DiodeTransistorPmos: -3.44399e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outVoltageBiasXXnXX0: 0.580001  V
** outVoltageBiasXXpXX1: 2.21601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21901  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.01701  V
** sourceGCC2: 3.01701  V


.END