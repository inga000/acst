** Name: two_stage_single_output_op_amp_51_8

.MACRO two_stage_single_output_op_amp_51_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=24e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=40e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=40e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=561e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=7e-6 W=599e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=8e-6 W=21e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=160e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=70e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=70e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=568e-6
mFoldedCascodeFirstStageLoad17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=160e-6
mMainBias18 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=115e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=46e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.5e-12
.EOM two_stage_single_output_op_amp_51_8

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 6.53301 mW
** Area: 10593 (mu_m)^2
** Transit frequency: 4.13701 MHz
** Transit frequency with error factor: 4.13664 MHz
** Slew rate: 3.89987 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 4.25 V
** VoutMin: 0.550001 V
** VcmMax: 5.12001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorPmos: -5.49679e+07 muA
** NormalTransistorPmos: -2.21509e+07 muA
** NormalTransistorPmos: -2.16599e+07 muA
** NormalTransistorPmos: -3.39699e+07 muA
** NormalTransistorPmos: -2.16599e+07 muA
** NormalTransistorPmos: -3.39699e+07 muA
** NormalTransistorNmos: 2.16591e+07 muA
** NormalTransistorNmos: 2.16591e+07 muA
** DiodeTransistorNmos: 2.16591e+07 muA
** NormalTransistorNmos: 2.46171e+07 muA
** NormalTransistorNmos: 1.23091e+07 muA
** NormalTransistorNmos: 1.23091e+07 muA
** NormalTransistorNmos: 1.14161e+09 muA
** NormalTransistorNmos: 1.14161e+09 muA
** NormalTransistorPmos: -1.1416e+09 muA
** DiodeTransistorNmos: 5.49671e+07 muA
** DiodeTransistorNmos: 2.21501e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** outVoltageBiasXXnXX1: 1.15501  V
** outVoltageBiasXXnXX2: 0.560001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.605001  V
** out1: 1.32101  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.92401  V
** innerStageBias: 0.355001  V


.END