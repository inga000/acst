.suckt  two_stage_single_output_op_amp_191_10 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m4 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
m5 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m6 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourceNmos sourceNmos nmos
m7 FirstStageYout1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m8 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m10 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c2 out sourceNmos 
m13 out ibias sourceNmos sourceNmos nmos
m14 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
m16 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m17 ibias ibias sourceNmos sourceNmos nmos
m18 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m19 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_191_10

