** Name: two_stage_single_output_op_amp_46_9

.MACRO two_stage_single_output_op_amp_46_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=11e-6
m2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=33e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=296e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=22e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
m6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=251e-6
m7 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=35e-6
m8 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=296e-6
m9 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=180e-6
m10 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=180e-6
m11 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=98e-6
m12 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=98e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
m14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=179e-6
m15 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=79e-6
m16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=235e-6
m17 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=35e-6
m18 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=251e-6
m19 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=541e-6
m20 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=541e-6
m21 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=293e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 17e-12
.EOM two_stage_single_output_op_amp_46_9

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 14.1321 mW
** Area: 14997 (mu_m)^2
** Transit frequency: 5.85101 MHz
** Transit frequency with error factor: 5.85111 MHz
** Slew rate: 5.92963 V/mu_s
** Phase margin: 60.1606°
** CMRR: 132 dB
** VoutMax: 4.25 V
** VoutMin: 1.62001 V
** VcmMax: 3.93001 V
** VcmMin: -0.279999 V


** Expected Currents: 
** NormalTransistorPmos: -8.52039e+07 muA
** NormalTransistorPmos: -3.79699e+07 muA
** NormalTransistorNmos: 1.01082e+08 muA
** NormalTransistorNmos: 1.72177e+08 muA
** NormalTransistorNmos: 1.01084e+08 muA
** NormalTransistorNmos: 1.72179e+08 muA
** DiodeTransistorPmos: -1.01081e+08 muA
** DiodeTransistorPmos: -1.01082e+08 muA
** NormalTransistorPmos: -1.01083e+08 muA
** NormalTransistorPmos: -1.01082e+08 muA
** NormalTransistorPmos: -1.4219e+08 muA
** NormalTransistorPmos: -7.10959e+07 muA
** NormalTransistorPmos: -7.10959e+07 muA
** NormalTransistorNmos: 2.33881e+09 muA
** DiodeTransistorNmos: 2.33881e+09 muA
** NormalTransistorPmos: -2.3388e+09 muA
** DiodeTransistorNmos: 8.52031e+07 muA
** NormalTransistorNmos: 8.52021e+07 muA
** DiodeTransistorNmos: 3.79691e+07 muA
** DiodeTransistorNmos: 3.79701e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.15201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.02601  V
** inputVoltageBiasXXnXX2: 1.33001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 1.01301  V
** outSourceVoltageBiasXXnXX2: 0.692001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.28601  V
** innerTransistorStack2Load2: 4.28701  V
** out1: 3.32201  V
** sourceGCC1: 0.762001  V
** sourceGCC2: 0.762001  V
** sourceTransconductance: 3.29001  V
** inner: 1.01301  V


.END