.suckt  two_stage_single_output_op_amp_7_9 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m3 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerOutputLoad1 sourceNmos sourceNmos nmos
m4 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerOutputLoad1 sourceNmos sourceNmos nmos
m6 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c2 out sourceNmos 
m9 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m10 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m11 out outFirstStage sourcePmos sourcePmos pmos
m12 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m14 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_7_9

