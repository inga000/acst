** Name: two_stage_single_output_op_amp_4_1

.MACRO two_stage_single_output_op_amp_4_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=10e-6 W=73e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=142e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=142e-6
mSecondStage1Transconductor5 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=174e-6
mSimpleFirstStageLoad6 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=10e-6 W=73e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=17e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=56e-6
mSecondStage1StageBias9 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=393e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=17e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_4_1

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 2.36001 mW
** Area: 6258 (mu_m)^2
** Transit frequency: 2.92201 MHz
** Transit frequency with error factor: 2.91578 MHz
** Slew rate: 12.58 V/mu_s
** Phase margin: 72.7657°
** CMRR: 90 dB
** negPSRR: 87 dB
** posPSRR: 93 dB
** VoutMax: 4.66001 V
** VoutMin: 0.370001 V
** VcmMax: 3.42001 V
** VcmMin: 0.610001 V


** Expected Currents: 
** DiodeTransistorNmos: 2.85291e+07 muA
** DiodeTransistorNmos: 2.85281e+07 muA
** NormalTransistorNmos: 2.85291e+07 muA
** NormalTransistorNmos: 2.85281e+07 muA
** NormalTransistorPmos: -5.70589e+07 muA
** NormalTransistorPmos: -2.85299e+07 muA
** NormalTransistorPmos: -2.85299e+07 muA
** NormalTransistorNmos: 3.94986e+08 muA
** NormalTransistorPmos: -3.94985e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.10001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.773001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 1.17801  V
** innerSourceLoad1: 0.559001  V
** innerTransistorStack2Load1: 0.558001  V
** sourceTransconductance: 3.74601  V


.END