.suckt  two_stage_single_output_op_amp_175_1 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mMainBias2 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad5 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad7 FirstStageYout1 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad8 outFirstStage ibias sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1Transconductor13 out outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias14 out inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mMainBias15 ibias ibias sourceNmos sourceNmos nmos
mMainBias16 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mMainBias17 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_175_1

