** Name: symmetrical_op_amp116

.MACRO symmetrical_op_amp116 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=9e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=26e-6
mMainBias3 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=340e-6
mSymmetricalFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=28e-6
mSecondStage1StageBias6 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=67e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias7 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=67e-6
mSymmetricalFirstStageTransconductor8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=20e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias9 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=4e-6 W=68e-6
mSecondStage1StageBias10 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=90e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=20e-6
mMainBias12 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=7e-6 W=32e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=140e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=19e-6
mSymmetricalFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=8e-6 W=19e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=56e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=8e-6 W=56e-6
mMainBias18 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=156e-6
mSymmetricalFirstStageLoad19 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=76e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor20 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=226e-6
mSecondStage1Transconductor21 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=226e-6
mSymmetricalFirstStageLoad22 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=76e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp116

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 1.94701 mW
** Area: 6013 (mu_m)^2
** Transit frequency: 2.50701 MHz
** Transit frequency with error factor: 2.50702 MHz
** Slew rate: 4.53322 V/mu_s
** Phase margin: 76.2034°
** CMRR: 139 dB
** negPSRR: 132 dB
** posPSRR: 60 dB
** VoutMax: 4.25 V
** VoutMin: 0.330001 V
** VcmMax: 4.81001 V
** VcmMin: 0.990001 V


** Expected Currents: 
** NormalTransistorNmos: 1.53208e+08 muA
** NormalTransistorNmos: 3.55351e+07 muA
** NormalTransistorPmos: -6.90439e+07 muA
** NormalTransistorPmos: -1.52889e+07 muA
** NormalTransistorPmos: -1.52899e+07 muA
** NormalTransistorPmos: -1.52889e+07 muA
** NormalTransistorPmos: -1.52899e+07 muA
** NormalTransistorNmos: 3.05761e+07 muA
** NormalTransistorNmos: 1.52881e+07 muA
** NormalTransistorNmos: 1.52881e+07 muA
** NormalTransistorNmos: 4.54871e+07 muA
** NormalTransistorNmos: 4.54861e+07 muA
** NormalTransistorPmos: -4.54879e+07 muA
** NormalTransistorPmos: -4.54869e+07 muA
** NormalTransistorNmos: 4.54871e+07 muA
** NormalTransistorNmos: 4.54861e+07 muA
** NormalTransistorPmos: -4.54879e+07 muA
** NormalTransistorPmos: -4.54869e+07 muA
** DiodeTransistorNmos: 6.90431e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.53207e+08 muA
** DiodeTransistorPmos: -3.55359e+07 muA


** Expected Voltages: 
** ibias: 0.707001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.761001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.584001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 4.27801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.80901  V
** innerStageBias: 0.201001  V
** innerTransconductance: 4.40001  V
** inner: 0.179001  V
** inner: 4.40001  V


.END