** Name: two_stage_single_output_op_amp_61_9

.MACRO two_stage_single_output_op_amp_61_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=29e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=7e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=550e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=45e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=9e-6 W=186e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=37e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=20e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=550e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=20e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=135e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=9e-6 W=353e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=45e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=52e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=52e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=24e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=9e-6 W=522e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=131e-6
mFoldedCascodeFirstStageLoad22 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=49e-6
mMainBias23 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=9e-6 W=155e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_61_9

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 4.78601 mW
** Area: 14770 (mu_m)^2
** Transit frequency: 3.82701 MHz
** Transit frequency with error factor: 3.82699 MHz
** Slew rate: 4.21646 V/mu_s
** Phase margin: 61.8795°
** CMRR: 142 dB
** VoutMax: 4.25 V
** VoutMin: 0.740001 V
** VcmMax: 3.24001 V
** VcmMin: -0.379999 V


** Expected Currents: 
** NormalTransistorNmos: 1.84928e+08 muA
** NormalTransistorPmos: -8.44799e+06 muA
** NormalTransistorPmos: -2.81969e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 2.85691e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 2.85691e+07 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90469e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -9.52299e+06 muA
** NormalTransistorPmos: -9.52299e+06 muA
** NormalTransistorNmos: 6.58465e+08 muA
** DiodeTransistorNmos: 6.58464e+08 muA
** NormalTransistorPmos: -6.58464e+08 muA
** DiodeTransistorNmos: 8.44701e+06 muA
** NormalTransistorNmos: 8.44601e+06 muA
** DiodeTransistorNmos: 2.81961e+07 muA
** DiodeTransistorNmos: 2.81971e+07 muA
** DiodeTransistorPmos: -1.84927e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.14001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.14601  V
** outSourceVoltageBiasXXnXX1: 0.573001  V
** outSourceVoltageBiasXXnXX2: 0.584001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.54701  V
** innerTransistorStack2Load2: 4.45801  V
** out1: 4.16901  V
** sourceGCC1: 0.585001  V
** sourceGCC2: 0.585001  V
** sourceTransconductance: 3.23901  V
** inner: 0.572001  V


.END