** Name: two_stage_single_output_op_amp_188_9

.MACRO two_stage_single_output_op_amp_188_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=23e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=9e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=79e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=336e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=29e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=128e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=79e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=23e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=336e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=6e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=128e-6
mSimpleFirstStageLoad15 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=186e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=444e-6
mSimpleFirstStageLoad17 outFirstStage ibias sourcePmos sourcePmos pmos4 L=5e-6 W=186e-6
mMainBias18 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=41e-6
mMainBias19 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=114e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.30001e-12
.EOM two_stage_single_output_op_amp_188_9

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 8.53601 mW
** Area: 10094 (mu_m)^2
** Transit frequency: 6.17501 MHz
** Transit frequency with error factor: 6.16219 MHz
** Slew rate: 5.82001 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 1.20001 V
** VcmMax: 5.09001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorPmos: -1.43189e+07 muA
** NormalTransistorPmos: -3.96289e+07 muA
** NormalTransistorNmos: 4.09381e+07 muA
** NormalTransistorNmos: 4.09391e+07 muA
** DiodeTransistorNmos: 4.09381e+07 muA
** NormalTransistorPmos: -6.53189e+07 muA
** NormalTransistorPmos: -6.53189e+07 muA
** NormalTransistorNmos: 4.87591e+07 muA
** DiodeTransistorNmos: 4.87581e+07 muA
** NormalTransistorNmos: 2.43801e+07 muA
** NormalTransistorNmos: 2.43801e+07 muA
** NormalTransistorNmos: 1.50271e+09 muA
** DiodeTransistorNmos: 1.50271e+09 muA
** NormalTransistorPmos: -1.5027e+09 muA
** DiodeTransistorNmos: 1.43181e+07 muA
** NormalTransistorNmos: 1.43171e+07 muA
** DiodeTransistorNmos: 3.96281e+07 muA
** NormalTransistorNmos: 3.96291e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.12401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.22801  V
** outInputVoltageBiasXXnXX2: 1.60401  V
** outSourceVoltageBiasXXnXX1: 0.614001  V
** outSourceVoltageBiasXXnXX2: 0.802001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.10301  V
** out1: 2.14601  V
** sourceTransconductance: 1.94501  V
** inner: 0.612001  V
** inner: 0.803001  V


.END