.suckt  symmetrical_op_amp20 ibias in1 in2 out sourceNmos sourcePmos
m1 outFirstStage outFirstStage sourcePmos sourcePmos pmos
m2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m3 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m4 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m5 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m6 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos
m7 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m8 out outFirstStage sourcePmos sourcePmos pmos
m9 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m10 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m11 ibias ibias sourceNmos sourceNmos nmos
.end symmetrical_op_amp20

