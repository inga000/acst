.suckt  two_stage_fully_differential_op_amp_31_7 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m5 outFeedback outFeedback sourceNmos sourceNmos nmos
m6 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m7 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m8 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m9 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m10 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m12 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m13 FirstStageYinnerTransistorStack1Load1 outFeedback sourceNmos sourceNmos nmos
m14 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m15 FirstStageYinnerTransistorStack2Load1 outFeedback sourceNmos sourceNmos nmos
m16 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m17 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m18 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m19 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m20 out1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m21 out1 out1FirstStage sourcePmos sourcePmos pmos
m22 out2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m23 out2 out2FirstStage sourcePmos sourcePmos pmos
m24 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m25 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m26 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m27 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m28 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_31_7

