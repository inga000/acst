** Name: two_stage_single_output_op_amp_71_9

.MACRO two_stage_single_output_op_amp_71_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=36e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=135e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=594e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=89e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=33e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=27e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=12e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=11e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=135e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=594e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=55e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=89e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=89e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=482e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=338e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=55e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=345e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.90001e-12
.EOM two_stage_single_output_op_amp_71_9

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 4.81501 mW
** Area: 9931 (mu_m)^2
** Transit frequency: 2.56601 MHz
** Transit frequency with error factor: 2.56228 MHz
** Slew rate: 3.77436 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** VoutMax: 4.25 V
** VoutMin: 0.700001 V
** VcmMax: 5.12001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorPmos: -1.28563e+08 muA
** NormalTransistorPmos: -1.81664e+08 muA
** NormalTransistorPmos: -2.23369e+07 muA
** NormalTransistorPmos: -3.35439e+07 muA
** NormalTransistorPmos: -2.23369e+07 muA
** NormalTransistorPmos: -3.35439e+07 muA
** DiodeTransistorNmos: 2.23361e+07 muA
** NormalTransistorNmos: 2.23361e+07 muA
** NormalTransistorNmos: 2.24111e+07 muA
** NormalTransistorNmos: 2.24101e+07 muA
** NormalTransistorNmos: 1.12061e+07 muA
** NormalTransistorNmos: 1.12061e+07 muA
** NormalTransistorNmos: 5.65675e+08 muA
** DiodeTransistorNmos: 5.65675e+08 muA
** NormalTransistorPmos: -5.65674e+08 muA
** DiodeTransistorNmos: 1.28564e+08 muA
** NormalTransistorNmos: 1.28564e+08 muA
** DiodeTransistorNmos: 1.81665e+08 muA
** DiodeTransistorNmos: 1.81664e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.20801  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.560001  V
** outSourceVoltageBiasXXpXX1: 4.14701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.648001  V
** out1: 0.567001  V
** sourceGCC1: 4.18601  V
** sourceGCC2: 4.18601  V
** sourceTransconductance: 1.85901  V
** inner: 0.555001  V


.END