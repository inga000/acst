.suckt  two_stage_single_output_op_amp_87_9 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mMainBias2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mMainBias3 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mMainBias4 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mTelescopicFirstStageLoad5 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mTelescopicFirstStageLoad6 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mTelescopicFirstStageLoad7 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
mTelescopicFirstStageLoad8 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mTelescopicFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos
mTelescopicFirstStageStageBias10 sourceTransconductance ibias sourcePmos sourcePmos pmos
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mSecondStage1StageBias14 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos
mMainBias16 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mMainBias17 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mMainBias18 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias19 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias20 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
mMainBias21 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_87_9

