.suckt  symmetrical_op_amp69 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mSymmetricalFirstStageLoad2 outFirstStage outFirstStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad3 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageStageBias4 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
mSymmetricalFirstStageStageBias5 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mSymmetricalFirstStageTransconductor6 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSymmetricalFirstStageTransconductor7 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1StageBias8 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos
mSecondStage1StageBias9 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStage1Transconductor10 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias12 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor13 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mMainBias15 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mMainBias16 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mSecondStage1StageBias17 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
.end symmetrical_op_amp69

