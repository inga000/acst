** Name: one_stage_single_output_op_amp110

.MACRO one_stage_single_output_op_amp110 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=33e-6
mTelescopicFirstStageLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=33e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=26e-6
mTelescopicFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=427e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=5e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=33e-6
mTelescopicFirstStageLoad8 out FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=33e-6
mMainBias9 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=68e-6
mTelescopicFirstStageLoad10 FirstStageYinnerOutputLoad2 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=30e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=84e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=84e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=26e-6
mMainBias14 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=7e-6
mTelescopicFirstStageLoad15 out outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=30e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=427e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp110

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 0.949001 mW
** Area: 3929 (mu_m)^2
** Transit frequency: 2.86301 MHz
** Transit frequency with error factor: 2.86283 MHz
** Slew rate: 8.34599 V/mu_s
** Phase margin: 88.8085°
** CMRR: 138 dB
** VoutMax: 3.07001 V
** VoutMin: 0.820001 V
** VcmMax: 3 V
** VcmMin: 1.15001 V


** Expected Currents: 
** NormalTransistorNmos: 3.75121e+07 muA
** NormalTransistorPmos: -2.73799e+06 muA
** NormalTransistorPmos: -6.47759e+07 muA
** NormalTransistorPmos: -6.47759e+07 muA
** DiodeTransistorNmos: 6.47751e+07 muA
** NormalTransistorNmos: 6.47741e+07 muA
** NormalTransistorNmos: 6.47751e+07 muA
** DiodeTransistorNmos: 6.47741e+07 muA
** NormalTransistorPmos: -1.67061e+08 muA
** DiodeTransistorPmos: -1.6706e+08 muA
** NormalTransistorPmos: -6.47749e+07 muA
** NormalTransistorPmos: -6.47749e+07 muA
** DiodeTransistorNmos: 2.73701e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -3.75129e+07 muA


** Expected Voltages: 
** ibias: 3.36001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.566001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.18101  V
** outVoltageBiasXXpXX2: 1.93801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.42201  V
** innerOutputLoad2: 1.22501  V
** innerSourceLoad2: 0.668001  V
** innerTransistorStack1Load2: 0.667001  V
** sourceGCC1: 2.99401  V
** sourceGCC2: 2.99401  V
** inner: 4.17701  V


.END