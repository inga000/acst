.suckt  symmetrical_op_amp171 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage out2FirstStage out1FirstStage out1FirstStage pmos
m2 out1FirstStage out1FirstStage sourcePmos sourcePmos pmos
m3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage pmos
m4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m5 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m7 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m8 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m9 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m10 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m11 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m12 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m13 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos
m14 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m15 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m17 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m18 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
.end symmetrical_op_amp171

