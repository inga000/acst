** Name: two_stage_single_output_op_amp_3_6

.MACRO two_stage_single_output_op_amp_3_6 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=177e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=30e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=36e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=116e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=177e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=295e-6
mSecondStage1Transconductor9 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=416e-6
mSimpleFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=119e-6
mMainBias11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=15e-6
mSimpleFirstStageTransconductor12 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=70e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=167e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=36e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=64e-6
mSecondStage1StageBias16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=116e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=70e-6
mMainBias18 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=83e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.9001e-12
.EOM two_stage_single_output_op_amp_3_6

** Expected Performance Values: 
** Gain: 132 dB
** Power consumption: 2.92601 mW
** Area: 7858 (mu_m)^2
** Transit frequency: 3.06201 MHz
** Transit frequency with error factor: 3.0542 MHz
** Slew rate: 5.86976 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** negPSRR: 94 dB
** posPSRR: 114 dB
** VoutMax: 3.23001 V
** VoutMin: 0.310001 V
** VcmMax: 3.47001 V
** VcmMin: 0.200001 V


** Expected Currents: 
** NormalTransistorNmos: 5.94611e+07 muA
** NormalTransistorPmos: -8.41509e+07 muA
** NormalTransistorPmos: -6.42909e+07 muA
** DiodeTransistorNmos: 8.46581e+07 muA
** NormalTransistorNmos: 8.46581e+07 muA
** NormalTransistorNmos: 8.46581e+07 muA
** NormalTransistorPmos: -1.69316e+08 muA
** NormalTransistorPmos: -8.46589e+07 muA
** NormalTransistorPmos: -8.46589e+07 muA
** NormalTransistorNmos: 1.87957e+08 muA
** NormalTransistorNmos: 1.87956e+08 muA
** NormalTransistorPmos: -1.87956e+08 muA
** DiodeTransistorPmos: -1.87957e+08 muA
** DiodeTransistorNmos: 8.41501e+07 muA
** DiodeTransistorNmos: 6.42901e+07 muA
** DiodeTransistorPmos: -5.94619e+07 muA
** NormalTransistorPmos: -5.94619e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.759001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.66201  V
** outSourceVoltageBiasXXpXX1: 3.83101  V
** outVoltageBiasXXnXX0: 0.712001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.79701  V
** innerTransconductance: 0.190001  V
** inner: 3.83101  V


.END