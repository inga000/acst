.suckt  one_stage_fully_differential_op_amp3 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
m1 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m3 outFeedback outFeedback sourceNmos sourceNmos nmos
m4 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m5 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m6 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m7 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m8 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m9 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m10 out1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m11 FirstStageYinnerTransistorStack1Load1 outFeedback sourceNmos sourceNmos nmos
m12 out2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m13 FirstStageYinnerTransistorStack2Load1 outFeedback sourceNmos sourceNmos nmos
m14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m15 out1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m16 out2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c1 out1 sourceNmos 
c2 out2 sourceNmos 
m17 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m18 ibias ibias sourcePmos sourcePmos pmos
.end one_stage_fully_differential_op_amp3

