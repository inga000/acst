** Name: two_stage_single_output_op_amp_62_1

.MACRO two_stage_single_output_op_amp_62_1 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=23e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=42e-6
m3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=7e-6
m4 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=9e-6 W=14e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=103e-6
m7 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=63e-6
m8 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=49e-6
m9 inputVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=28e-6
m10 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=180e-6
m11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=8e-6 W=33e-6
m12 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=11e-6
m13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=8e-6 W=33e-6
m14 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=118e-6
m15 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=118e-6
m16 out inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=590e-6
m17 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=176e-6
m18 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=63e-6
m19 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=78e-6
m20 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=78e-6
m21 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=9e-6 W=103e-6
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=14e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_62_1

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 3.72001 mW
** Area: 11084 (mu_m)^2
** Transit frequency: 3.60301 MHz
** Transit frequency with error factor: 3.60309 MHz
** Slew rate: 4.09624 V/mu_s
** Phase margin: 61.3065°
** CMRR: 136 dB
** VoutMax: 4.65001 V
** VoutMin: 0.550001 V
** VcmMax: 3.08001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.61901e+06 muA
** NormalTransistorNmos: 1.16661e+07 muA
** NormalTransistorNmos: 6.73301e+06 muA
** NormalTransistorNmos: 1.86091e+07 muA
** NormalTransistorNmos: 2.80941e+07 muA
** NormalTransistorNmos: 1.86091e+07 muA
** NormalTransistorNmos: 2.80941e+07 muA
** DiodeTransistorPmos: -1.86099e+07 muA
** NormalTransistorPmos: -1.86099e+07 muA
** NormalTransistorPmos: -1.86099e+07 muA
** NormalTransistorPmos: -1.89729e+07 muA
** DiodeTransistorPmos: -1.89739e+07 muA
** NormalTransistorPmos: -9.48599e+06 muA
** NormalTransistorPmos: -9.48599e+06 muA
** NormalTransistorNmos: 6.56688e+08 muA
** NormalTransistorPmos: -6.56687e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.61999e+06 muA
** NormalTransistorPmos: -2.62099e+06 muA
** DiodeTransistorPmos: -1.16669e+07 muA
** DiodeTransistorPmos: -6.73399e+06 muA


** Expected Voltages: 
** ibias: 1.16201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.68601  V
** inputVoltageBiasXXpXX3: 4.08201  V
** out: 2.5  V
** outFirstStage: 0.957001  V
** outInputVoltageBiasXXpXX1: 3.26001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.13001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.43801  V
** out1: 4.07401  V
** sourceGCC1: 0.525001  V
** sourceGCC2: 0.525001  V
** sourceTransconductance: 3.24801  V
** inner: 4.13001  V


.END