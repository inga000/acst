** Name: two_stage_single_output_op_amp_187_10

.MACRO two_stage_single_output_op_amp_187_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=18e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
m3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=57e-6
m5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m6 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=31e-6
m7 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=70e-6
m8 out ibias sourceNmos sourceNmos nmos4 L=8e-6 W=315e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=9e-6 W=48e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=5e-6
m11 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=69e-6
m12 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
m13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=5e-6
m14 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=140e-6
m15 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=285e-6
m16 outFirstStage inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=498e-6
m17 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=40e-6
m18 FirstStageYout1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=498e-6
m19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=388e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_187_10

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 2.71801 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 3.07401 MHz
** Transit frequency with error factor: 3.03942 MHz
** Slew rate: 6.96629 V/mu_s
** Phase margin: 60.1606°
** CMRR: 86 dB
** VoutMax: 4.66001 V
** VoutMin: 0.230001 V
** VcmMax: 5.04001 V
** VcmMin: 1.61001 V


** Expected Currents: 
** NormalTransistorNmos: 3.88921e+07 muA
** NormalTransistorNmos: 1.71331e+07 muA
** NormalTransistorPmos: -1.20229e+07 muA
** NormalTransistorNmos: 1.27942e+08 muA
** NormalTransistorNmos: 1.27943e+08 muA
** DiodeTransistorNmos: 1.27942e+08 muA
** NormalTransistorPmos: -1.46987e+08 muA
** NormalTransistorPmos: -1.46987e+08 muA
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorNmos: 3.80921e+07 muA
** NormalTransistorNmos: 1.90461e+07 muA
** NormalTransistorNmos: 1.90461e+07 muA
** NormalTransistorNmos: 1.71554e+08 muA
** NormalTransistorPmos: -1.71553e+08 muA
** NormalTransistorPmos: -1.71554e+08 muA
** DiodeTransistorNmos: 1.20221e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.88929e+07 muA
** DiodeTransistorPmos: -1.71339e+07 muA


** Expected Voltages: 
** ibias: 0.633001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.96801  V
** inputVoltageBiasXXpXX2: 4.07101  V
** out: 2.5  V
** outFirstStage: 4.27801  V
** outVoltageBiasXXnXX1: 0.783001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.228001  V
** out1: 2.09501  V
** sourceTransconductance: 1.66901  V
** innerTransconductance: 4.71501  V


.END