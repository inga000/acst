** Name: two_stage_single_output_op_amp_62_5

.MACRO two_stage_single_output_op_amp_62_5 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=15e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m3 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=10e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=128e-6
m5 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=2e-6 W=8e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=175e-6
m7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=442e-6
m8 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
m9 inputVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=26e-6
m10 out outFirstStage sourceNmos sourceNmos nmos4 L=10e-6 W=334e-6
m11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=39e-6
m12 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=53e-6
m13 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=30e-6
m14 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=39e-6
m15 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=107e-6
m16 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=107e-6
m17 out outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=442e-6
m18 outFirstStage inputVoltageBiasXXpXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=8e-6 W=184e-6
m19 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
m20 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=126e-6
m21 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=126e-6
m22 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=175e-6
m23 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
m24 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=128e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 7.20001e-12
.EOM two_stage_single_output_op_amp_62_5

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 4.70701 mW
** Area: 11694 (mu_m)^2
** Transit frequency: 5.00201 MHz
** Transit frequency with error factor: 5.00166 MHz
** Slew rate: 4.64709 V/mu_s
** Phase margin: 60.1606°
** CMRR: 142 dB
** VoutMax: 3.55001 V
** VoutMin: 0.530001 V
** VcmMax: 3.30001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.52371e+07 muA
** NormalTransistorNmos: 1.42851e+07 muA
** NormalTransistorNmos: 1.25051e+07 muA
** NormalTransistorNmos: 3.36751e+07 muA
** NormalTransistorNmos: 5.09491e+07 muA
** NormalTransistorNmos: 3.36751e+07 muA
** NormalTransistorNmos: 5.09491e+07 muA
** DiodeTransistorPmos: -3.36759e+07 muA
** NormalTransistorPmos: -3.36759e+07 muA
** NormalTransistorPmos: -3.36759e+07 muA
** NormalTransistorPmos: -3.45509e+07 muA
** DiodeTransistorPmos: -3.45519e+07 muA
** NormalTransistorPmos: -1.72749e+07 muA
** NormalTransistorPmos: -1.72749e+07 muA
** NormalTransistorNmos: 7.77453e+08 muA
** NormalTransistorPmos: -7.77452e+08 muA
** DiodeTransistorPmos: -7.77453e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.52379e+07 muA
** NormalTransistorPmos: -2.52389e+07 muA
** DiodeTransistorPmos: -1.42859e+07 muA
** NormalTransistorPmos: -1.42869e+07 muA
** DiodeTransistorPmos: -1.25059e+07 muA


** Expected Voltages: 
** ibias: 1.13701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX3: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.932001  V
** outInputVoltageBiasXXpXX1: 3.45001  V
** outInputVoltageBiasXXpXX2: 2.98201  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.22501  V
** outSourceVoltageBiasXXpXX2: 3.99101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.53501  V
** out1: 4.21001  V
** sourceGCC1: 0.529001  V
** sourceGCC2: 0.529001  V
** sourceTransconductance: 3.21501  V
** inner: 4.22401  V
** inner: 3.99101  V


.END