** Name: two_stage_single_output_op_amp_60_1

.MACRO two_stage_single_output_op_amp_60_1 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=17e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
m3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=119e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=97e-6
m5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=8e-6
m6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=66e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=221e-6
m8 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=21e-6
m9 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=73e-6
m10 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=56e-6
m11 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=21e-6
m12 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=88e-6
m13 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=88e-6
m14 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=460e-6
m15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=37e-6
m16 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=66e-6
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=59e-6
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=59e-6
m19 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=97e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=119e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_60_1

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 4.78101 mW
** Area: 10781 (mu_m)^2
** Transit frequency: 2.65301 MHz
** Transit frequency with error factor: 2.65287 MHz
** Slew rate: 3.53688 V/mu_s
** Phase margin: 73.9116°
** CMRR: 138 dB
** VoutMax: 4.35001 V
** VoutMin: 0.570001 V
** VcmMax: 3.18001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.00571e+07 muA
** NormalTransistorNmos: 1.52981e+07 muA
** NormalTransistorNmos: 1.59681e+07 muA
** NormalTransistorNmos: 2.40241e+07 muA
** NormalTransistorNmos: 1.59681e+07 muA
** NormalTransistorNmos: 2.40241e+07 muA
** NormalTransistorPmos: -1.59689e+07 muA
** NormalTransistorPmos: -1.59689e+07 muA
** DiodeTransistorPmos: -1.59689e+07 muA
** NormalTransistorPmos: -1.61149e+07 muA
** DiodeTransistorPmos: -1.61159e+07 muA
** NormalTransistorPmos: -8.05699e+06 muA
** NormalTransistorPmos: -8.05699e+06 muA
** NormalTransistorNmos: 8.62726e+08 muA
** NormalTransistorPmos: -8.62725e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.00579e+07 muA
** NormalTransistorPmos: -2.00589e+07 muA
** DiodeTransistorPmos: -1.52989e+07 muA


** Expected Voltages: 
** ibias: 1.18101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.976001  V
** outInputVoltageBiasXXpXX1: 3.39801  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXpXX2: 3.78501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.08601  V
** out1: 3.30201  V
** sourceGCC1: 0.524001  V
** sourceGCC2: 0.524001  V
** sourceTransconductance: 3.27801  V
** inner: 4.19901  V


.END