** Name: two_stage_single_output_op_amp_106_3

.MACRO two_stage_single_output_op_amp_106_3 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=194e-6
m2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=93e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=93e-6
m4 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos4 L=8e-6 W=59e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=28e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=354e-6
m7 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
m8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=6e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=101e-6
m10 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=93e-6
m11 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=43e-6
m12 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=330e-6
m13 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=93e-6
m14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=8e-6 W=600e-6
m15 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=42e-6
m16 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=6e-6
m17 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=354e-6
m18 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=6e-6
m19 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=36e-6
m20 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=36e-6
m21 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=152e-6
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.5e-12
.EOM two_stage_single_output_op_amp_106_3

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 2.13501 mW
** Area: 14815 (mu_m)^2
** Transit frequency: 2.53301 MHz
** Transit frequency with error factor: 2.53332 MHz
** Slew rate: 7.25395 V/mu_s
** Phase margin: 60.1606°
** CMRR: 124 dB
** VoutMax: 3.31001 V
** VoutMin: 0.300001 V
** VcmMax: 3 V
** VcmMin: 1.46001 V


** Expected Currents: 
** NormalTransistorNmos: 1.17481e+07 muA
** NormalTransistorNmos: 9.00071e+07 muA
** NormalTransistorPmos: -5.27869e+07 muA
** NormalTransistorPmos: -2.95229e+07 muA
** NormalTransistorPmos: -2.95229e+07 muA
** DiodeTransistorNmos: 2.95221e+07 muA
** DiodeTransistorNmos: 2.95221e+07 muA
** NormalTransistorNmos: 2.95221e+07 muA
** NormalTransistorNmos: 2.95221e+07 muA
** NormalTransistorPmos: -1.49056e+08 muA
** DiodeTransistorPmos: -1.49057e+08 muA
** NormalTransistorPmos: -2.95239e+07 muA
** NormalTransistorPmos: -2.95239e+07 muA
** NormalTransistorNmos: 1.9343e+08 muA
** NormalTransistorPmos: -1.93429e+08 muA
** NormalTransistorPmos: -1.93428e+08 muA
** DiodeTransistorNmos: 5.27861e+07 muA
** DiodeTransistorPmos: -1.17489e+07 muA
** NormalTransistorPmos: -1.175e+07 muA
** DiodeTransistorPmos: -9.00079e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.84501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outInputVoltageBiasXXpXX1: 3.56401  V
** outSourceVoltageBiasXXpXX1: 4.28201  V
** outSourceVoltageBiasXXpXX3: 3.68501  V
** outVoltageBiasXXpXX2: 1.48501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.62801  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 2.96201  V
** sourceGCC2: 2.95401  V
** innerStageBias: 3.78701  V
** inner: 4.28101  V


.END