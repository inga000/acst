** Name: two_stage_single_output_op_amp_73_5

.MACRO two_stage_single_output_op_amp_73_5 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=15e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=105e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=9e-6 W=23e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=8e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=562e-6
m7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=23e-6
m8 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=134e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=84e-6
m10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=8e-6 W=84e-6
m11 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=135e-6
m12 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=111e-6
m13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=105e-6
m14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=28e-6
m15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=28e-6
m16 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=57e-6
m17 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=562e-6
m18 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=9e-6 W=28e-6
m19 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=9e-6 W=28e-6
m20 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=28e-6
m21 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=28e-6
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 5.60001e-12
.EOM two_stage_single_output_op_amp_73_5

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 9.54701 mW
** Area: 11878 (mu_m)^2
** Transit frequency: 4.01301 MHz
** Transit frequency with error factor: 4.01326 MHz
** Slew rate: 3.54627 V/mu_s
** Phase margin: 60.1606°
** CMRR: 137 dB
** VoutMax: 3.24001 V
** VoutMin: 0.5 V
** VcmMax: 4.66001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorNmos: 2.57131e+07 muA
** NormalTransistorNmos: 2.56711e+07 muA
** NormalTransistorPmos: -2e+07 muA
** NormalTransistorPmos: -3.06669e+07 muA
** NormalTransistorPmos: -2e+07 muA
** NormalTransistorPmos: -3.06669e+07 muA
** NormalTransistorNmos: 1.99991e+07 muA
** NormalTransistorNmos: 1.99991e+07 muA
** DiodeTransistorNmos: 1.99991e+07 muA
** NormalTransistorNmos: 2.13311e+07 muA
** NormalTransistorNmos: 2.13301e+07 muA
** NormalTransistorNmos: 1.06661e+07 muA
** NormalTransistorNmos: 1.06661e+07 muA
** NormalTransistorNmos: 1.78672e+09 muA
** NormalTransistorPmos: -1.78671e+09 muA
** DiodeTransistorPmos: -1.78671e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.57139e+07 muA
** NormalTransistorPmos: -2.57149e+07 muA
** DiodeTransistorPmos: -2.56719e+07 muA
** DiodeTransistorPmos: -2.56709e+07 muA


** Expected Voltages: 
** ibias: 1.24001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.37601  V
** out: 2.5  V
** outFirstStage: 0.905001  V
** outInputVoltageBiasXXpXX1: 2.67401  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.83701  V
** outSourceVoltageBiasXXpXX2: 3.69001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerStageBias: 0.624001  V
** out1: 1.11001  V
** sourceGCC1: 3.53701  V
** sourceGCC2: 3.53701  V
** sourceTransconductance: 1.94501  V
** inner: 3.83501  V


.END