** Name: symmetrical_op_amp79

.MACRO symmetrical_op_amp79 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=10e-6
m2 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=8e-6 W=108e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
m4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=16e-6
m5 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=8e-6
m6 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=314e-6
m7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=6e-6
m8 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=314e-6
m9 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=27e-6
m10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=183e-6
m11 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
m12 out outVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=558e-6
m13 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=183e-6
m14 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=600e-6
m15 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=8e-6 W=108e-6
m16 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
m17 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=3e-6 W=239e-6
m18 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=239e-6
m19 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=90e-6
m20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=371e-6
m21 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=371e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp79

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 7.70501 mW
** Area: 12207 (mu_m)^2
** Transit frequency: 23.1541 MHz
** Transit frequency with error factor: 23.1541 MHz
** Slew rate: 35.4107 V/mu_s
** Phase margin: 60.7336°
** CMRR: 141 dB
** negPSRR: 49 dB
** posPSRR: 42 dB
** VoutMax: 4.27001 V
** VoutMin: 0.730001 V
** VcmMax: 4.61001 V
** VcmMin: 1.43001 V


** Expected Currents: 
** NormalTransistorNmos: 1.20881e+07 muA
** NormalTransistorNmos: 2.70741e+07 muA
** NormalTransistorPmos: -1.79144e+08 muA
** DiodeTransistorPmos: -2.99003e+08 muA
** DiodeTransistorPmos: -2.99003e+08 muA
** NormalTransistorNmos: 5.98006e+08 muA
** DiodeTransistorNmos: 5.98005e+08 muA
** NormalTransistorNmos: 2.99004e+08 muA
** NormalTransistorNmos: 2.99004e+08 muA
** NormalTransistorNmos: 3.57345e+08 muA
** NormalTransistorNmos: 3.57344e+08 muA
** NormalTransistorPmos: -3.57344e+08 muA
** NormalTransistorPmos: -3.57343e+08 muA
** DiodeTransistorNmos: 3.57345e+08 muA
** NormalTransistorPmos: -3.57344e+08 muA
** NormalTransistorPmos: -3.57343e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 1.79145e+08 muA
** DiodeTransistorPmos: -1.20889e+07 muA
** DiodeTransistorPmos: -2.70749e+07 muA


** Expected Voltages: 
** ibias: 1.18501  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 4.20501  V
** innerComplementarySecondStage: 0.962001  V
** inputVoltageBiasXXpXX0: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.20501  V
** outSourceVoltageBiasXXnXX1: 0.593001  V
** outVoltageBiasXXnXX2: 1.13601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.85401  V
** innerStageBias: 0.557001  V
** innerTransconductance: 4.74901  V
** inner: 4.74901  V
** inner: 0.591001  V


.END