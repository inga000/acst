** Name: one_stage_single_output_op_amp55

.MACRO one_stage_single_output_op_amp55 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=61e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=61e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=15e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=158e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=61e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=54e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=54e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=119e-6
mMainBias10 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=89e-6
mFoldedCascodeFirstStageLoad11 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=3e-6 W=61e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=254e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=256e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=256e-6
mFoldedCascodeFirstStageLoad15 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=254e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp55

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 2.36401 mW
** Area: 2991 (mu_m)^2
** Transit frequency: 5.28801 MHz
** Transit frequency with error factor: 5.28832 MHz
** Slew rate: 5.13835 V/mu_s
** Phase margin: 88.2356°
** CMRR: 140 dB
** VoutMax: 4.09001 V
** VoutMin: 0.850001 V
** VcmMax: 5.21001 V
** VcmMin: 0.870001 V


** Expected Currents: 
** NormalTransistorNmos: 1.10555e+08 muA
** NormalTransistorPmos: -1.03157e+08 muA
** NormalTransistorPmos: -1.7617e+08 muA
** NormalTransistorPmos: -1.03157e+08 muA
** NormalTransistorPmos: -1.7617e+08 muA
** DiodeTransistorNmos: 1.03158e+08 muA
** NormalTransistorNmos: 1.03157e+08 muA
** NormalTransistorNmos: 1.03158e+08 muA
** DiodeTransistorNmos: 1.03157e+08 muA
** NormalTransistorNmos: 1.46025e+08 muA
** NormalTransistorNmos: 7.30121e+07 muA
** NormalTransistorNmos: 7.30121e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.10554e+08 muA
** DiodeTransistorPmos: -1.10555e+08 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.23901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.604001  V
** innerTransistorStack1Load2: 0.602001  V
** out1: 1.25301  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.87601  V


.END