.suckt  symmetrical_op_amp111 ibias in1 in2 out sourceNmos sourcePmos
mSymmetricalFirstStageLoad1 out2FirstStage out2FirstStage out1FirstStage out1FirstStage pmos
mSymmetricalFirstStageLoad2 out1FirstStage out1FirstStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage pmos
mSymmetricalFirstStageLoad4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSymmetricalFirstStageTransconductor6 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSymmetricalFirstStageTransconductor7 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1StageBias8 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos
mSecondStage1StageBias9 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStage1Transconductor10 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor11 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias12 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor13 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mMainBias15 ibias ibias sourceNmos sourceNmos nmos
.end symmetrical_op_amp111

