** Name: two_stage_single_output_op_amp_79_8

.MACRO two_stage_single_output_op_amp_79_8 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=90e-6
m3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m5 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=281e-6
m6 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=11e-6
m7 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
m8 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=93e-6
m9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=93e-6
m10 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=11e-6
m11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=15e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=15e-6
m13 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=15e-6
m14 SecondStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=342e-6
m15 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=535e-6
m16 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=55e-6
m17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=280e-6
m18 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=204e-6
m19 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=55e-6
m20 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
m21 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.80001e-12
.EOM two_stage_single_output_op_amp_79_8

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 6.83001 mW
** Area: 7167 (mu_m)^2
** Transit frequency: 3.97101 MHz
** Transit frequency with error factor: 3.97111 MHz
** Slew rate: 3.58863 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 4.25 V
** VoutMin: 0.340001 V
** VcmMax: 5.17001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorPmos: -2.83885e+08 muA
** NormalTransistorPmos: -2.02879e+08 muA
** NormalTransistorPmos: -2.44699e+07 muA
** NormalTransistorPmos: -4.15689e+07 muA
** NormalTransistorPmos: -2.44699e+07 muA
** NormalTransistorPmos: -4.15689e+07 muA
** NormalTransistorNmos: 2.44691e+07 muA
** NormalTransistorNmos: 2.44681e+07 muA
** NormalTransistorNmos: 2.44691e+07 muA
** NormalTransistorNmos: 2.44681e+07 muA
** NormalTransistorNmos: 3.41951e+07 muA
** NormalTransistorNmos: 3.41941e+07 muA
** NormalTransistorNmos: 1.70981e+07 muA
** NormalTransistorNmos: 1.70981e+07 muA
** NormalTransistorNmos: 7.7601e+08 muA
** NormalTransistorNmos: 7.76009e+08 muA
** NormalTransistorPmos: -7.76009e+08 muA
** DiodeTransistorNmos: 2.83886e+08 muA
** DiodeTransistorNmos: 2.0288e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.955001  V
** outVoltageBiasXXnXX2: 0.569001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.386001  V
** innerTransistorStack1Load2: 0.388001  V
** innerTransistorStack2Load2: 0.388001  V
** out1: 0.581001  V
** sourceGCC1: 4.11901  V
** sourceGCC2: 4.11901  V
** sourceTransconductance: 1.89401  V
** innerStageBias: 0.369001  V


.END