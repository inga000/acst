.suckt  two_stage_fully_differential_op_amp_30_3 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_2 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_Load_3 outFeedback outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_4 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m_FullyDifferential_FeedbackdStage_StageBias_5 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_6 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackStage_Transconductor_8 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_9 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_10 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FeedbackStage_Transconductor_11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FirstStage_Load_12 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m_FullyDifferential_FirstStage_Load_13 FirstStageYinnerTransistorStack1Load1 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_14 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m_FullyDifferential_FirstStage_Load_15 FirstStageYinnerTransistorStack2Load1 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_StageBias_16 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m_FullyDifferential_FirstStage_StageBias_17 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Transconductor_18 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_FullyDifferential_FirstStage_Transconductor_19 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_Transconductor_20 out1 out1FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_21 out1 ibias SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m_FullyDifferential_SecondStage1_StageBias_22 SecondStage1YinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_Transconductor_23 out2 out2FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_StageBias_24 out2 ibias SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m_FullyDifferential_SecondStage2_StageBias_25 SecondStage2YinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_26 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_27 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_FullyDifferential_MainBias_28 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_30_3

