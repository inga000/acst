** Name: two_stage_single_output_op_amp_44_8

.MACRO two_stage_single_output_op_amp_44_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=13e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=72e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=112e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=423e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=318e-6
mFoldedCascodeFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad11 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=72e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=50e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=50e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=7e-6 W=254e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=290e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=362e-6
mFoldedCascodeFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=9e-6 W=275e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_44_8

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 5.12801 mW
** Area: 10537 (mu_m)^2
** Transit frequency: 4.96501 MHz
** Transit frequency with error factor: 4.96534 MHz
** Slew rate: 4.1539 V/mu_s
** Phase margin: 64.1713°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.75 V
** VcmMax: 4.09001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorPmos: -2.57479e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 3.04981e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 3.04981e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -2.29029e+07 muA
** NormalTransistorPmos: -1.14519e+07 muA
** NormalTransistorPmos: -1.14519e+07 muA
** NormalTransistorNmos: 9.18883e+08 muA
** NormalTransistorNmos: 9.18882e+08 muA
** NormalTransistorPmos: -9.18882e+08 muA
** DiodeTransistorNmos: 2.57471e+07 muA
** DiodeTransistorNmos: 2.57481e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.12301  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.565001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.11301  V
** out1: 3.36201  V
** sourceGCC1: 0.568001  V
** sourceGCC2: 0.568001  V
** sourceTransconductance: 3.22401  V
** innerStageBias: 0.533001  V


.END