.suckt  symmetrical_op_amp26 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos
mSymmetricalFirstStageLoad2 outFirstStage outFirstStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad3 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSymmetricalFirstStageTransconductor5 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSymmetricalFirstStageTransconductor6 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1StageBias7 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
mSecondStage1StageBias8 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStage1Transconductor9 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias11 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos
mSecondStageWithVoltageBiasAsStageBiasStageBias12 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor13 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mMainBias15 ibias ibias sourceNmos sourceNmos nmos
mSecondStage1StageBias16 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
.end symmetrical_op_amp26

