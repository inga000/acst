** Name: two_stage_single_output_op_amp_71_1

.MACRO two_stage_single_output_op_amp_71_1 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=24e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=15e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=60e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=110e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=35e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=22e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=22e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=13e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=75e-6
mFoldedCascodeFirstStageLoad11 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=24e-6
mMainBias12 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=426e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=207e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=125e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mSecondStage1StageBias17 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=378e-6
mFoldedCascodeFirstStageLoad18 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=125e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_71_1

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 3.54201 mW
** Area: 4973 (mu_m)^2
** Transit frequency: 3.92701 MHz
** Transit frequency with error factor: 3.9237 MHz
** Slew rate: 3.70067 V/mu_s
** Phase margin: 63.0254°
** CMRR: 106 dB
** VoutMax: 4.78001 V
** VoutMin: 0.230001 V
** VcmMax: 5.18001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 2.03068e+08 muA
** NormalTransistorNmos: 9.95591e+07 muA
** NormalTransistorPmos: -1.67629e+07 muA
** NormalTransistorPmos: -2.51429e+07 muA
** NormalTransistorPmos: -1.67649e+07 muA
** NormalTransistorPmos: -2.51469e+07 muA
** DiodeTransistorNmos: 1.67641e+07 muA
** NormalTransistorNmos: 1.67641e+07 muA
** NormalTransistorNmos: 1.67611e+07 muA
** NormalTransistorNmos: 1.67601e+07 muA
** NormalTransistorNmos: 8.38101e+06 muA
** NormalTransistorNmos: 8.38101e+06 muA
** NormalTransistorNmos: 3.45418e+08 muA
** NormalTransistorPmos: -3.45417e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.03067e+08 muA
** DiodeTransistorPmos: -9.95599e+07 muA


** Expected Voltages: 
** ibias: 1.13701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.638001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.21101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.484001  V
** out1: 0.645001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V


.END