** Name: two_stage_single_output_op_amp_195_9

.MACRO two_stage_single_output_op_amp_195_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=9e-6 W=13e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=12e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=143e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=35e-6
mMainBias7 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=41e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=87e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=10e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=13e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=34e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=143e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=9e-6 W=13e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=13e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=309e-6
mMainBias17 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=80e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=209e-6
mSimpleFirstStageLoad19 outFirstStage ibias sourcePmos sourcePmos pmos4 L=2e-6 W=309e-6
mMainBias20 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=597e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.80001e-12
.EOM two_stage_single_output_op_amp_195_9

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 12.2921 mW
** Area: 4803 (mu_m)^2
** Transit frequency: 5.31801 MHz
** Transit frequency with error factor: 5.31046 MHz
** Slew rate: 5.01248 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 1.24001 V
** VcmMax: 5.24001 V
** VcmMin: 1.52001 V


** Expected Currents: 
** NormalTransistorPmos: -1.45739e+08 muA
** NormalTransistorPmos: -1.96489e+07 muA
** DiodeTransistorNmos: 5.07191e+07 muA
** DiodeTransistorNmos: 5.07201e+07 muA
** NormalTransistorNmos: 5.07191e+07 muA
** NormalTransistorNmos: 5.07201e+07 muA
** NormalTransistorPmos: -7.54809e+07 muA
** NormalTransistorPmos: -7.54809e+07 muA
** NormalTransistorNmos: 4.95211e+07 muA
** NormalTransistorNmos: 4.95201e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.12207e+09 muA
** DiodeTransistorNmos: 2.12207e+09 muA
** NormalTransistorPmos: -2.12206e+09 muA
** DiodeTransistorNmos: 1.4574e+08 muA
** NormalTransistorNmos: 1.45741e+08 muA
** DiodeTransistorNmos: 1.96481e+07 muA
** DiodeTransistorNmos: 1.96471e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.39301  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.64401  V
** outSourceVoltageBiasXXnXX1: 0.822001  V
** outSourceVoltageBiasXXnXX2: 0.621001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.14301  V
** innerStageBias: 0.640001  V
** innerTransistorStack2Load1: 1.14301  V
** out1: 2.19501  V
** sourceTransconductance: 1.94501  V
** inner: 0.823001  V


.END