** Name: two_stage_single_output_op_amp_206_7

.MACRO two_stage_single_output_op_amp_206_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=7e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=11e-6
m3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
m4 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=30e-6
m5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
m6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=42e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=9e-6
m8 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=89e-6
m9 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=30e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=7e-6
m11 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=7e-6
m12 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
m13 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=11e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
m15 out outFirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=556e-6
m16 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=388e-6
m17 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=9e-6
m18 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=31e-6
m19 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=388e-6
m20 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=166e-6
m21 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=166e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_206_7

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 5.34301 mW
** Area: 11284 (mu_m)^2
** Transit frequency: 2.75 MHz
** Transit frequency with error factor: 2.74825 MHz
** Slew rate: 3.50005 V/mu_s
** Phase margin: 67.6091°
** CMRR: 121 dB
** VoutMax: 4.25 V
** VoutMin: 0.640001 V
** VcmMax: 4.58001 V
** VcmMin: 1.71001 V


** Expected Currents: 
** NormalTransistorPmos: -1.01939e+07 muA
** NormalTransistorPmos: -3.51119e+07 muA
** DiodeTransistorNmos: 1.79917e+08 muA
** NormalTransistorNmos: 1.79918e+08 muA
** NormalTransistorNmos: 1.79919e+08 muA
** DiodeTransistorNmos: 1.79918e+08 muA
** NormalTransistorPmos: -1.88017e+08 muA
** NormalTransistorPmos: -1.88018e+08 muA
** NormalTransistorPmos: -1.88019e+08 muA
** NormalTransistorPmos: -1.88018e+08 muA
** NormalTransistorNmos: 1.62031e+07 muA
** DiodeTransistorNmos: 1.62021e+07 muA
** NormalTransistorNmos: 8.10101e+06 muA
** NormalTransistorNmos: 8.10101e+06 muA
** NormalTransistorNmos: 6.27255e+08 muA
** NormalTransistorPmos: -6.27254e+08 muA
** DiodeTransistorNmos: 1.01931e+07 muA
** NormalTransistorNmos: 1.01921e+07 muA
** DiodeTransistorNmos: 3.51111e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.14001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.50601  V
** outSourceVoltageBiasXXnXX1: 0.753001  V
** outSourceVoltageBiasXXpXX1: 3.93501  V
** outVoltageBiasXXnXX2: 1.04701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack1Load1: 1.15601  V
** innerTransistorStack1Load2: 4.03201  V
** innerTransistorStack2Load2: 4.03201  V
** sourceTransconductance: 1.89201  V
** inner: 0.753001  V


.END