** Name: one_stage_single_output_op_amp116

.MACRO one_stage_single_output_op_amp116 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=6e-6
mTelescopicFirstStageStageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=59e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=43e-6
mTelescopicFirstStageLoad4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=16e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=9e-6
mTelescopicFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=92e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=53e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=53e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias10 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mTelescopicFirstStageLoad11 out outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=92e-6
mTelescopicFirstStageStageBias12 sourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=59e-6
mTelescopicFirstStageLoad13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=16e-6
mTelescopicFirstStageLoad14 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=113e-6
mMainBias15 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=42e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp116

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 0.585001 mW
** Area: 3226 (mu_m)^2
** Transit frequency: 2.66901 MHz
** Transit frequency with error factor: 2.66905 MHz
** Slew rate: 4.8308 V/mu_s
** Phase margin: 81.933°
** CMRR: 150 dB
** VoutMax: 3.43001 V
** VoutMin: 1.10001 V
** VcmMax: 3.69001 V
** VcmMin: 1.35001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00561e+07 muA
** NormalTransistorPmos: -4.64549e+07 muA
** NormalTransistorNmos: 2.52371e+07 muA
** NormalTransistorNmos: 2.52361e+07 muA
** NormalTransistorPmos: -2.52379e+07 muA
** NormalTransistorPmos: -2.52369e+07 muA
** DiodeTransistorPmos: -2.52379e+07 muA
** NormalTransistorNmos: 9.69291e+07 muA
** DiodeTransistorNmos: 9.69301e+07 muA
** NormalTransistorNmos: 2.52371e+07 muA
** NormalTransistorNmos: 2.52371e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 4.64541e+07 muA
** DiodeTransistorPmos: -1.00569e+07 muA


** Expected Voltages: 
** ibias: 1.20501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.68601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.603001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 3.59201  V
** out1: 2.87001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.601001  V


.END