** Name: two_stage_single_output_op_amp_65_1

.MACRO two_stage_single_output_op_amp_65_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=11e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=66e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=14e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=14e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=66e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=66e-6
mMainBias8 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=215e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=166e-6
mFoldedCascodeFirstStageLoad10 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=14e-6
mMainBias11 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=33e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=67e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=67e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=7e-6 W=153e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=7e-6 W=211e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=586e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=153e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_65_1

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 3.38301 mW
** Area: 9338 (mu_m)^2
** Transit frequency: 3.44501 MHz
** Transit frequency with error factor: 3.44519 MHz
** Slew rate: 3.69204 V/mu_s
** Phase margin: 63.0254°
** CMRR: 142 dB
** VoutMax: 4.68001 V
** VoutMin: 0.580001 V
** VcmMax: 3.21001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 8.18991e+07 muA
** NormalTransistorNmos: 1.26161e+07 muA
** NormalTransistorNmos: 1.67301e+07 muA
** NormalTransistorNmos: 2.51421e+07 muA
** NormalTransistorNmos: 1.67301e+07 muA
** NormalTransistorNmos: 2.51421e+07 muA
** NormalTransistorPmos: -1.67309e+07 muA
** NormalTransistorPmos: -1.67319e+07 muA
** NormalTransistorPmos: -1.67309e+07 muA
** NormalTransistorPmos: -1.67319e+07 muA
** NormalTransistorPmos: -1.68269e+07 muA
** NormalTransistorPmos: -1.68279e+07 muA
** NormalTransistorPmos: -8.41299e+06 muA
** NormalTransistorPmos: -8.41299e+06 muA
** NormalTransistorNmos: 5.21825e+08 muA
** NormalTransistorPmos: -5.21824e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -8.18999e+07 muA
** DiodeTransistorPmos: -1.26169e+07 muA


** Expected Voltages: 
** ibias: 1.19101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.73601  V
** out: 2.5  V
** outFirstStage: 0.986001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX2: 4.12001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.47601  V
** innerTransistorStack1Load2: 4.50601  V
** innerTransistorStack2Load2: 4.50601  V
** out1: 4.26801  V
** sourceGCC1: 0.519001  V
** sourceGCC2: 0.519001  V
** sourceTransconductance: 3.23501  V


.END