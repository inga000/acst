** Name: two_stage_single_output_op_amp_78_5

.MACRO two_stage_single_output_op_amp_78_5 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=3e-6 W=26e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=30e-6
mMainBias3 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=39e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=95e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=8e-6 W=14e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=12e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=480e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=18e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=3e-6 W=26e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=49e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=49e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=95e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=39e-6
mMainBias14 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=69e-6
mSecondStage1Transconductor15 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=590e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=30e-6
mMainBias17 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=215e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=8e-6 W=28e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=32e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=32e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=480e-6
mFoldedCascodeFirstStageLoad23 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=8e-6 W=28e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.40001e-12
.EOM two_stage_single_output_op_amp_78_5

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 11.6731 mW
** Area: 11828 (mu_m)^2
** Transit frequency: 4.64301 MHz
** Transit frequency with error factor: 4.64257 MHz
** Slew rate: 3.51596 V/mu_s
** Phase margin: 60.1606°
** CMRR: 137 dB
** VoutMax: 3.42001 V
** VoutMin: 0.510001 V
** VcmMax: 4.74001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 5.45741e+07 muA
** NormalTransistorNmos: 1.77671e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -3.10909e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -3.10909e+07 muA
** DiodeTransistorNmos: 1.90471e+07 muA
** DiodeTransistorNmos: 1.90461e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90461e+07 muA
** NormalTransistorNmos: 2.40851e+07 muA
** DiodeTransistorNmos: 2.40861e+07 muA
** NormalTransistorNmos: 1.20421e+07 muA
** NormalTransistorNmos: 1.20421e+07 muA
** NormalTransistorNmos: 2.19008e+09 muA
** NormalTransistorPmos: -2.19007e+09 muA
** DiodeTransistorPmos: -2.19007e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.45749e+07 muA
** NormalTransistorPmos: -5.45759e+07 muA
** DiodeTransistorPmos: -1.77679e+07 muA
** DiodeTransistorPmos: -1.77689e+07 muA


** Expected Voltages: 
** ibias: 1.13901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.46001  V
** out: 2.5  V
** outFirstStage: 0.916001  V
** outInputVoltageBiasXXpXX1: 2.85801  V
** outSourceVoltageBiasXXnXX1: 0.570001  V
** outSourceVoltageBiasXXpXX1: 3.92901  V
** outSourceVoltageBiasXXpXX2: 3.77401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.566001  V
** innerTransistorStack2Load2: 0.566001  V
** out1: 1.12101  V
** sourceGCC1: 3.57401  V
** sourceGCC2: 3.57401  V
** sourceTransconductance: 1.94201  V
** inner: 0.569001  V
** inner: 3.92401  V


.END