.suckt  symmetrical_op_amp18 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mMainBias2 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad4 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSymmetricalFirstStageTransconductor6 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSymmetricalFirstStageTransconductor7 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1StageBias8 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
mSecondStage1StageBias9 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStage1Transconductor10 out outFirstStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias11 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos
mSecondStageWithVoltageBiasAsStageBiasStageBias12 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor13 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mMainBias14 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
mMainBias15 ibias ibias sourceNmos sourceNmos nmos
mMainBias16 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end symmetrical_op_amp18

