.suckt  two_stage_fully_differential_op_amp_45_6 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 outVoltageBiasXXpXX3 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m4 outVoltageBiasXXpXX4 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m5 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m6 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m7 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m8 outFeedback outFeedback sourceNmos sourceNmos nmos
m9 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m10 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m11 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m15 out1FirstStage outVoltageBiasXXpXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m16 out2FirstStage outVoltageBiasXXpXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m17 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m18 FirstStageYinnerTransistorStack1Load2 outFeedback sourceNmos sourceNmos nmos
m19 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m20 FirstStageYinnerTransistorStack2Load2 outFeedback sourceNmos sourceNmos nmos
m21 sourceTransconductance outVoltageBiasXXpXX4 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m22 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
m23 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m24 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m25 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m26 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m27 out1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m28 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m29 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m30 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m31 out2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m32 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m33 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m34 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m35 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m36 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m37 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m38 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m39 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourceTransconductance sourceTransconductance pmos
m40 outVoltageBiasXXpXX4 outVoltageBiasXXpXX4 sourcePmos sourcePmos pmos
m41 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_45_6

