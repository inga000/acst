** Name: one_stage_single_output_op_amp116

.MACRO one_stage_single_output_op_amp116 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=10e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=235e-6
m3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=24e-6
m4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=14e-6
m5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=16e-6
m6 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=49e-6
m7 out outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=13e-6
m8 sourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=235e-6
m9 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=13e-6
m10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=26e-6
m11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=26e-6
m12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
m13 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=55e-6
m14 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=53e-6
m15 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=16e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp116

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 1.45501 mW
** Area: 3122 (mu_m)^2
** Transit frequency: 2.625 MHz
** Transit frequency with error factor: 2.62468 MHz
** Slew rate: 11.5822 V/mu_s
** Phase margin: 89.9544°
** CMRR: 143 dB
** VoutMax: 3.39001 V
** VoutMin: 1.14001 V
** VcmMax: 3.65001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorNmos: 4.90801e+07 muA
** NormalTransistorPmos: -1.8234e+08 muA
** NormalTransistorNmos: 2.47621e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorPmos: -2.47629e+07 muA
** NormalTransistorPmos: -2.47619e+07 muA
** DiodeTransistorPmos: -2.47629e+07 muA
** NormalTransistorNmos: 2.31864e+08 muA
** DiodeTransistorNmos: 2.31865e+08 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 1.82341e+08 muA
** DiodeTransistorPmos: -4.90809e+07 muA


** Expected Voltages: 
** ibias: 1.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.27001  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.622001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 3.54901  V
** out1: 2.82601  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.619001  V


.END