** Name: two_stage_single_output_op_amp_29_10

.MACRO two_stage_single_output_op_amp_29_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=10e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=219e-6
mMainBias4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=20e-6
mSecondStage1StageBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=362e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=37e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=372e-6
mMainBias9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
mMainBias10 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=237e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=6e-6 W=522e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=37e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSecondStage1Transconductor14 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=219e-6
mMainBias16 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=162e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.7001e-12
.EOM two_stage_single_output_op_amp_29_10

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 6.27501 mW
** Area: 11693 (mu_m)^2
** Transit frequency: 6.97201 MHz
** Transit frequency with error factor: 6.93214 MHz
** Slew rate: 16.7646 V/mu_s
** Phase margin: 60.1606°
** CMRR: 86 dB
** negPSRR: 116 dB
** posPSRR: 84 dB
** VoutMax: 4.56001 V
** VoutMin: 0.260001 V
** VcmMax: 4.63001 V
** VcmMin: 1.97001 V


** Expected Currents: 
** NormalTransistorNmos: 1.50111e+07 muA
** NormalTransistorNmos: 2.33528e+08 muA
** NormalTransistorPmos: -1.22694e+08 muA
** DiodeTransistorPmos: -1.77565e+08 muA
** NormalTransistorPmos: -1.77565e+08 muA
** NormalTransistorNmos: 3.5513e+08 muA
** NormalTransistorNmos: 3.55129e+08 muA
** NormalTransistorNmos: 1.77566e+08 muA
** NormalTransistorNmos: 1.77566e+08 muA
** NormalTransistorNmos: 5.18693e+08 muA
** NormalTransistorPmos: -5.18692e+08 muA
** NormalTransistorPmos: -5.18693e+08 muA
** DiodeTransistorNmos: 1.22695e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.50119e+07 muA
** DiodeTransistorPmos: -2.33527e+08 muA


** Expected Voltages: 
** ibias: 0.670001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.81901  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.21701  V
** outVoltageBiasXXnXX1: 0.820001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.265001  V
** out1: 4.22201  V
** sourceTransconductance: 1.34501  V
** innerTransconductance: 4.46901  V


.END