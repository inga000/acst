** Name: two_stage_single_output_op_amp_8_10

.MACRO two_stage_single_output_op_amp_8_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
m2 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
m3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=143e-6
m4 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=32e-6
m5 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=591e-6
m6 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=200e-6
m7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=32e-6
m8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=143e-6
m9 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=143e-6
m10 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
m11 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=550e-6
Capacitor1 outFirstStage out 11.6001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_8_10

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 3.15601 mW
** Area: 5723 (mu_m)^2
** Transit frequency: 5.62701 MHz
** Transit frequency with error factor: 5.61691 MHz
** Slew rate: 8.0603 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** negPSRR: 152 dB
** posPSRR: 95 dB
** VoutMax: 4.61001 V
** VoutMin: 0.180001 V
** VcmMax: 4.65001 V
** VcmMin: 0.810001 V


** Expected Currents: 
** NormalTransistorNmos: 1.31994e+08 muA
** DiodeTransistorPmos: -4.69359e+07 muA
** NormalTransistorPmos: -4.69359e+07 muA
** NormalTransistorNmos: 9.38711e+07 muA
** NormalTransistorNmos: 4.69351e+07 muA
** NormalTransistorNmos: 4.69351e+07 muA
** NormalTransistorNmos: 3.95255e+08 muA
** NormalTransistorPmos: -3.95254e+08 muA
** NormalTransistorPmos: -3.95255e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.31993e+08 muA


** Expected Voltages: 
** ibias: 0.582001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.23601  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.24401  V
** sourceTransconductance: 1.86601  V
** innerTransconductance: 4.44201  V


.END