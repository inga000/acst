** Name: two_stage_single_output_op_amp_206_9

.MACRO two_stage_single_output_op_amp_206_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=30e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=9e-6
mMainBias4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=5e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=128e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=42e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=9e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=30e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=27e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=8e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=9e-6
mMainBias13 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=128e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=30e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=27e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=167e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=167e-6
mSimpleFirstStageLoad19 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=390e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=596e-6
mSimpleFirstStageLoad21 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=390e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=16e-6
mMainBias23 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=23e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_206_9

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 5.56301 mW
** Area: 12742 (mu_m)^2
** Transit frequency: 2.95701 MHz
** Transit frequency with error factor: 2.95466 MHz
** Slew rate: 3.50007 V/mu_s
** Phase margin: 67.0361°
** CMRR: 122 dB
** VoutMax: 4.25 V
** VoutMin: 1.40001 V
** VcmMax: 4.58001 V
** VcmMin: 1.81001 V


** Expected Currents: 
** NormalTransistorPmos: -1.81219e+07 muA
** NormalTransistorPmos: -2.60509e+07 muA
** DiodeTransistorNmos: 1.79917e+08 muA
** NormalTransistorNmos: 1.79918e+08 muA
** NormalTransistorNmos: 1.79919e+08 muA
** DiodeTransistorNmos: 1.79918e+08 muA
** NormalTransistorPmos: -1.88027e+08 muA
** NormalTransistorPmos: -1.88028e+08 muA
** NormalTransistorPmos: -1.88029e+08 muA
** NormalTransistorPmos: -1.88028e+08 muA
** NormalTransistorNmos: 1.62231e+07 muA
** DiodeTransistorNmos: 1.62221e+07 muA
** NormalTransistorNmos: 8.11101e+06 muA
** NormalTransistorNmos: 8.11101e+06 muA
** NormalTransistorNmos: 6.72381e+08 muA
** DiodeTransistorNmos: 6.7238e+08 muA
** NormalTransistorPmos: -6.7238e+08 muA
** DiodeTransistorNmos: 1.81211e+07 muA
** NormalTransistorNmos: 1.81201e+07 muA
** DiodeTransistorNmos: 2.60501e+07 muA
** NormalTransistorNmos: 2.60491e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.14001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.62601  V
** outInputVoltageBiasXXnXX2: 1.80201  V
** outSourceVoltageBiasXXnXX1: 0.813001  V
** outSourceVoltageBiasXXnXX2: 0.901001  V
** outSourceVoltageBiasXXpXX1: 3.93501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack1Load1: 1.15601  V
** innerTransistorStack1Load2: 4.03101  V
** innerTransistorStack2Load2: 4.03101  V
** out1: 2.09501  V
** sourceTransconductance: 1.90601  V
** inner: 0.811001  V
** inner: 0.899001  V


.END