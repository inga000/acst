.suckt  two_stage_fully_differential_op_amp_39_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m4 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m5 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m6 outFeedback outFeedback sourceNmos sourceNmos nmos
m7 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m8 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m9 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m11 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m13 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m14 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m15 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m16 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m17 out1FirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m18 FirstStageYinnerTransistorStack1Load2 ibias sourcePmos sourcePmos pmos
m19 out2FirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m20 FirstStageYinnerTransistorStack2Load2 ibias sourcePmos sourcePmos pmos
m21 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m22 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m23 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m24 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m25 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m26 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m27 out1 outVoltageBiasXXpXX2 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m28 SecondStage1YinnerStageBias ibias sourcePmos sourcePmos pmos
m29 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m30 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m31 out2 outVoltageBiasXXpXX2 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m32 SecondStage2YinnerStageBias ibias sourcePmos sourcePmos pmos
m33 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m34 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m35 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m36 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m37 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m38 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_39_4

