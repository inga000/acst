** Name: two_stage_single_output_op_amp_6_5

.MACRO two_stage_single_output_op_amp_6_5 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=37e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=9e-6 W=37e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=10e-6 W=242e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=44e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=275e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=37e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=155e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=9e-6 W=37e-6
mMainBias10 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=40e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=10e-6 W=511e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=275e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mMainBias16 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=10e-6 W=256e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_6_5

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 1.62101 mW
** Area: 12964 (mu_m)^2
** Transit frequency: 3.07401 MHz
** Transit frequency with error factor: 3.07004 MHz
** Slew rate: 4.71573 V/mu_s
** Phase margin: 63.5984°
** CMRR: 101 dB
** negPSRR: 97 dB
** posPSRR: 102 dB
** VoutMax: 4 V
** VoutMin: 0.330001 V
** VcmMax: 4.04001 V
** VcmMin: 0.570001 V


** Expected Currents: 
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorPmos: -1.04769e+07 muA
** DiodeTransistorNmos: 1.06541e+07 muA
** NormalTransistorNmos: 1.06531e+07 muA
** NormalTransistorNmos: 1.06541e+07 muA
** DiodeTransistorNmos: 1.06531e+07 muA
** NormalTransistorPmos: -2.13099e+07 muA
** NormalTransistorPmos: -1.06549e+07 muA
** NormalTransistorPmos: -1.06549e+07 muA
** NormalTransistorNmos: 2.34358e+08 muA
** NormalTransistorPmos: -2.34357e+08 muA
** DiodeTransistorPmos: -2.34358e+08 muA
** DiodeTransistorNmos: 1.04761e+07 muA
** DiodeTransistorPmos: -3.80919e+07 muA
** NormalTransistorPmos: -3.80909e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.734001  V
** outInputVoltageBiasXXpXX1: 3.43401  V
** outSourceVoltageBiasXXpXX1: 4.21701  V
** outVoltageBiasXXnXX0: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.559001  V
** innerTransistorStack1Load1: 0.559001  V
** out1: 1.13901  V
** sourceTransconductance: 3.30701  V
** inner: 4.21801  V


.END