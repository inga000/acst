** Name: two_stage_single_output_op_amp_77_9

.MACRO two_stage_single_output_op_amp_77_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=29e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=82e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=308e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=376e-6
m5 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=82e-6
m6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=7e-6 W=12e-6
m7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
m8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m9 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=308e-6
m10 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=12e-6
m11 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=86e-6
m12 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=82e-6
m13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=56e-6
m14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=56e-6
m15 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=5e-6
m16 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=82e-6
m17 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=551e-6
m18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=178e-6
m19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=96e-6
m20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=298e-6
m21 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=96e-6
m22 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=59e-6
m23 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=59e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_77_9

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 8.69301 mW
** Area: 8762 (mu_m)^2
** Transit frequency: 6.41401 MHz
** Transit frequency with error factor: 6.41364 MHz
** Slew rate: 7.9063 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 4.25 V
** VoutMin: 0.820001 V
** VcmMax: 5.17001 V
** VcmMin: 1.80001 V


** Expected Currents: 
** NormalTransistorPmos: -3.00433e+08 muA
** NormalTransistorPmos: -1.79635e+08 muA
** NormalTransistorPmos: -3.89889e+07 muA
** NormalTransistorPmos: -5.98179e+07 muA
** NormalTransistorPmos: -3.89889e+07 muA
** NormalTransistorPmos: -5.98179e+07 muA
** DiodeTransistorNmos: 3.89881e+07 muA
** DiodeTransistorNmos: 3.89871e+07 muA
** NormalTransistorNmos: 3.89881e+07 muA
** NormalTransistorNmos: 3.89871e+07 muA
** NormalTransistorNmos: 4.16551e+07 muA
** NormalTransistorNmos: 4.16541e+07 muA
** NormalTransistorNmos: 2.08281e+07 muA
** NormalTransistorNmos: 2.08281e+07 muA
** NormalTransistorNmos: 1.11891e+09 muA
** DiodeTransistorNmos: 1.11891e+09 muA
** NormalTransistorPmos: -1.1189e+09 muA
** DiodeTransistorNmos: 3.00434e+08 muA
** NormalTransistorNmos: 3.00433e+08 muA
** DiodeTransistorNmos: 1.79636e+08 muA
** DiodeTransistorNmos: 1.79635e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.22401  V
** outSourceVoltageBiasXXnXX1: 0.612001  V
** outSourceVoltageBiasXXnXX2: 0.556001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.465001  V
** innerTransistorStack1Load2: 0.603001  V
** innerTransistorStack2Load2: 0.599001  V
** out1: 1.52401  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.88501  V
** inner: 0.610001  V


.END