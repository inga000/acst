** Name: two_stage_single_output_op_amp_89_2

.MACRO two_stage_single_output_op_amp_89_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=175e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=68e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=14e-6
mTelescopicFirstStageLoad5 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mTelescopicFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=6e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=367e-6
mMainBias9 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=56e-6
mSecondStage1Transconductor10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=92e-6
mTelescopicFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=6e-6
mTelescopicFirstStageLoad12 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=14e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=28e-6
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=28e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=255e-6
mSecondStage1StageBias16 out ibias sourcePmos sourcePmos pmos4 L=5e-6 W=591e-6
mTelescopicFirstStageLoad17 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=14e-6
mMainBias18 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=532e-6
mTelescopicFirstStageStageBias19 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=5e-6 W=242e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_89_2

** Expected Performance Values: 
** Gain: 155 dB
** Power consumption: 1.30001 mW
** Area: 13933 (mu_m)^2
** Transit frequency: 2.67201 MHz
** Transit frequency with error factor: 2.67189 MHz
** Slew rate: 3.56903 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.80001 V
** VoutMin: 0.300001 V
** VcmMax: 4.08001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 2.45701e+07 muA
** NormalTransistorPmos: -7.82909e+07 muA
** NormalTransistorPmos: -3.77169e+07 muA
** NormalTransistorPmos: -5.71499e+06 muA
** NormalTransistorPmos: -5.71499e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorPmos: -3.60019e+07 muA
** NormalTransistorPmos: -5.71599e+06 muA
** NormalTransistorPmos: -5.71599e+06 muA
** NormalTransistorNmos: 8.79211e+07 muA
** NormalTransistorNmos: 8.79201e+07 muA
** NormalTransistorPmos: -8.79219e+07 muA
** DiodeTransistorNmos: 7.82901e+07 muA
** DiodeTransistorNmos: 3.77161e+07 muA
** DiodeTransistorPmos: -2.45709e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.23301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXpXX1: 2.33701  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.622001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21501  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.05201  V
** sourceGCC2: 3.05201  V
** innerTransconductance: 0.150001  V


.END