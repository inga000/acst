** Name: two_stage_single_output_op_amp_108_3

.MACRO two_stage_single_output_op_amp_108_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=229e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=30e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos4 L=4e-6 W=11e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=52e-6
mTelescopicFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=333e-6
mMainBias6 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=9e-6 W=38e-6
mTelescopicFirstStageLoad8 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=195e-6
mTelescopicFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=156e-6
mTelescopicFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=156e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=429e-6
mTelescopicFirstStageLoad12 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=195e-6
mMainBias13 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=97e-6
mMainBias14 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=319e-6
mTelescopicFirstStageLoad15 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=9e-6 W=42e-6
mTelescopicFirstStageTransconductor16 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=117e-6
mTelescopicFirstStageTransconductor17 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=117e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=4e-6 W=293e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
mSecondStage1StageBias20 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=4e-6 W=600e-6
mTelescopicFirstStageLoad21 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=9e-6 W=42e-6
mMainBias22 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=4e-6 W=45e-6
mMainBias23 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=4e-6 W=18e-6
mTelescopicFirstStageStageBias24 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=333e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.8001e-12
.EOM two_stage_single_output_op_amp_108_3

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 6.40501 mW
** Area: 14566 (mu_m)^2
** Transit frequency: 3.53301 MHz
** Transit frequency with error factor: 3.53258 MHz
** Slew rate: 19.3323 V/mu_s
** Phase margin: 60.1606°
** CMRR: 128 dB
** VoutMax: 3.16001 V
** VoutMin: 0.290001 V
** VcmMax: 3 V
** VcmMin: 0.530001 V


** Expected Currents: 
** NormalTransistorNmos: 4.79411e+07 muA
** NormalTransistorNmos: 1.58441e+08 muA
** NormalTransistorPmos: -1.14529e+08 muA
** NormalTransistorPmos: -4.58119e+07 muA
** NormalTransistorPmos: -7.42819e+07 muA
** NormalTransistorPmos: -7.42819e+07 muA
** NormalTransistorNmos: 7.42811e+07 muA
** NormalTransistorNmos: 7.42811e+07 muA
** NormalTransistorNmos: 7.42811e+07 muA
** NormalTransistorNmos: 7.42811e+07 muA
** NormalTransistorPmos: -3.07007e+08 muA
** DiodeTransistorPmos: -3.07007e+08 muA
** NormalTransistorPmos: -7.42829e+07 muA
** NormalTransistorPmos: -7.42829e+07 muA
** NormalTransistorNmos: 7.45722e+08 muA
** NormalTransistorPmos: -7.45721e+08 muA
** NormalTransistorPmos: -7.4572e+08 muA
** DiodeTransistorNmos: 1.1453e+08 muA
** DiodeTransistorNmos: 4.58111e+07 muA
** DiodeTransistorPmos: -4.79419e+07 muA
** NormalTransistorPmos: -4.79409e+07 muA
** DiodeTransistorPmos: -1.5844e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.66801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.691001  V
** outInputVoltageBiasXXpXX1: 3.42001  V
** outSourceVoltageBiasXXpXX1: 4.21001  V
** outSourceVoltageBiasXXpXX3: 3.68501  V
** outVoltageBiasXXnXX0: 0.558001  V
** outVoltageBiasXXnXX1: 0.705001  V
** outVoltageBiasXXpXX2: 1.46401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.48401  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 2.96801  V
** sourceGCC2: 2.96801  V
** innerStageBias: 3.75701  V
** inner: 4.21101  V


.END