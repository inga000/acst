.suckt  two_stage_single_output_op_amp_179_2 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_6 outFirstStage FirstStageYinnerSourceLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_SingleOutput_FirstStage_Load_7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_8 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_9 outFirstStage inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_StageBias_10 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m_SingleOutput_FirstStage_StageBias_11 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Transconductor_12 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_SingleOutput_FirstStage_Transconductor_13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_Transconductor_14 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_SingleOutput_SecondStage1_Transconductor_15 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_16 out ibias sourcePmos sourcePmos pmos
m_SingleOutput_SecondStage1_StageBias_17 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_18 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_19 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_20 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_179_2

