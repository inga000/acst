** Name: two_stage_single_output_op_amp_169_1

.MACRO two_stage_single_output_op_amp_169_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=43e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=47e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=4e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=14e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=42e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=118e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=118e-6
mSimpleFirstStageLoad9 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=109e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=193e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=38e-6
mSimpleFirstStageLoad12 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=109e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=102e-6
mSimpleFirstStageStageBias14 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=45e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSimpleFirstStageTransconductor16 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=77e-6
mSimpleFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=3e-6 W=148e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=591e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=4e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=77e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_169_1

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 2.11601 mW
** Area: 14995 (mu_m)^2
** Transit frequency: 3.74601 MHz
** Transit frequency with error factor: 3.743 MHz
** Slew rate: 4.79845 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** VoutMax: 4.49001 V
** VoutMin: 0.310001 V
** VcmMax: 3 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 4.12561e+07 muA
** NormalTransistorNmos: 2.17371e+07 muA
** DiodeTransistorPmos: -1.35369e+07 muA
** DiodeTransistorPmos: -1.35369e+07 muA
** NormalTransistorPmos: -1.35369e+07 muA
** NormalTransistorPmos: -1.35369e+07 muA
** NormalTransistorNmos: 2.49711e+07 muA
** NormalTransistorNmos: 2.49721e+07 muA
** NormalTransistorNmos: 2.49711e+07 muA
** NormalTransistorNmos: 2.49721e+07 muA
** NormalTransistorPmos: -2.28709e+07 muA
** NormalTransistorPmos: -2.28719e+07 muA
** NormalTransistorPmos: -1.14349e+07 muA
** NormalTransistorPmos: -1.14349e+07 muA
** NormalTransistorNmos: 3.00171e+08 muA
** NormalTransistorPmos: -3.0017e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -4.12569e+07 muA
** DiodeTransistorPmos: -2.17379e+07 muA


** Expected Voltages: 
** ibias: 1.11701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.73001  V
** out: 2.5  V
** outFirstStage: 0.712001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX2: 3.92801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.68601  V
** innerStageBias: 4.45501  V
** innerTransistorStack1Load2: 0.556001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.556001  V
** out1: 2.37201  V
** sourceTransconductance: 3.26701  V


.END