.suckt  two_stage_fully_differential_op_amp_17_7 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m3 outFeedback outFeedback sourcePmos sourcePmos pmos
m4 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m5 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m6 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m7 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m8 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m9 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m10 out1FirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m11 FirstStageYsourceGCC1 outFeedback sourcePmos sourcePmos pmos
m12 out2FirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m13 FirstStageYsourceGCC2 outFeedback sourcePmos sourcePmos pmos
m14 out1FirstStage ibias sourceNmos sourceNmos nmos
m15 out2FirstStage ibias sourceNmos sourceNmos nmos
m16 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m19 out1 ibias sourceNmos sourceNmos nmos
m20 out1 out1FirstStage sourcePmos sourcePmos pmos
m21 out2 ibias sourceNmos sourceNmos nmos
m22 out2 out2FirstStage sourcePmos sourcePmos pmos
m23 ibias ibias sourceNmos sourceNmos nmos
m24 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_17_7

