** Name: two_stage_single_output_op_amp_36_7

.MACRO two_stage_single_output_op_amp_36_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=20e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=182e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=54e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=391e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=15e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=10e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mMainBias10 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=52e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=575e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=15e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=182e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=141e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=54e-6
mMainBias16 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=594e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_36_7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 4.68601 mW
** Area: 6828 (mu_m)^2
** Transit frequency: 4.58401 MHz
** Transit frequency with error factor: 4.57635 MHz
** Slew rate: 10.5617 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** negPSRR: 92 dB
** posPSRR: 86 dB
** VoutMax: 4.25 V
** VoutMin: 0.210001 V
** VcmMax: 3.85001 V
** VcmMin: 1.66001 V


** Expected Currents: 
** NormalTransistorNmos: 6.48261e+07 muA
** NormalTransistorPmos: -9.76839e+07 muA
** DiodeTransistorPmos: -2.43919e+07 muA
** DiodeTransistorPmos: -2.43929e+07 muA
** NormalTransistorPmos: -2.43939e+07 muA
** NormalTransistorPmos: -2.43929e+07 muA
** NormalTransistorNmos: 4.87851e+07 muA
** DiodeTransistorNmos: 4.87841e+07 muA
** NormalTransistorNmos: 2.43931e+07 muA
** NormalTransistorNmos: 2.43931e+07 muA
** NormalTransistorNmos: 7.15815e+08 muA
** NormalTransistorPmos: -7.15814e+08 muA
** DiodeTransistorNmos: 9.76831e+07 muA
** NormalTransistorNmos: 9.76821e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.48269e+07 muA


** Expected Voltages: 
** ibias: 0.615001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.27001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.28801  V
** outSourceVoltageBiasXXnXX1: 0.644001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.28601  V
** innerTransistorStack2Load1: 4.28701  V
** out1: 3.44801  V
** sourceTransconductance: 1.72701  V
** inner: 0.642001  V


.END