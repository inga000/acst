.suckt  complementary_op_amp10 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 FirstStageYinnerSourceLoadNmos outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m5 FirstStageYinnerTransistorStack1LoadPmos ibias sourcePmos sourcePmos pmos
m6 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m7 FirstStageYinnerTransistorStack2LoadPmos ibias sourcePmos sourcePmos pmos
m8 FirstStageYinnerSourceLoadNmos outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m9 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m10 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m11 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m12 FirstStageYsourceTransconductanceNmos inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m13 FirstStageYsourceTransconductancePmos ibias sourcePmos sourcePmos pmos
m14 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m15 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m16 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m17 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c1 out sourceNmos 
m18 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m19 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m20 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m21 ibias ibias sourcePmos sourcePmos pmos
.end complementary_op_amp10

