** Name: two_stage_single_output_op_amp_11_9

.MACRO two_stage_single_output_op_amp_11_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=28e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=352e-6
mSimpleFirstStageLoad4 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=10e-6 W=31e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=10e-6 W=77e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=8e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=28e-6
mSecondStage1StageBias10 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=352e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=8e-6
mMainBias12 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=10e-6 W=77e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=93e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=10e-6 W=31e-6
mMainBias16 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=113e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_11_9

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 2.66501 mW
** Area: 6541 (mu_m)^2
** Transit frequency: 3.03801 MHz
** Transit frequency with error factor: 3.03571 MHz
** Slew rate: 3.64187 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 100 dB
** posPSRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 0.960001 V
** VcmMax: 3.65001 V
** VcmMin: 0.790001 V


** Expected Currents: 
** NormalTransistorNmos: 5.58601e+06 muA
** NormalTransistorPmos: -3.70069e+07 muA
** DiodeTransistorPmos: -8.21499e+06 muA
** DiodeTransistorPmos: -8.21599e+06 muA
** NormalTransistorPmos: -8.21499e+06 muA
** NormalTransistorPmos: -8.21599e+06 muA
** NormalTransistorNmos: 1.64291e+07 muA
** NormalTransistorNmos: 8.21401e+06 muA
** NormalTransistorNmos: 8.21401e+06 muA
** NormalTransistorNmos: 4.63954e+08 muA
** DiodeTransistorNmos: 4.63953e+08 muA
** NormalTransistorPmos: -4.63953e+08 muA
** DiodeTransistorNmos: 3.70061e+07 muA
** NormalTransistorNmos: 3.70051e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.58699e+06 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.36601  V
** outSourceVoltageBiasXXnXX1: 0.683001  V
** outVoltageBiasXXpXX0: 4.24401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.24101  V
** innerTransistorStack1Load1: 4.19101  V
** innerTransistorStack2Load1: 4.18901  V
** sourceTransconductance: 1.90401  V
** inner: 0.681001  V


.END