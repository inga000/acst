** Name: two_stage_single_output_op_amp_78_3

.MACRO two_stage_single_output_op_amp_78_3 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=18e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=153e-6
m3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=5e-6 W=183e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=99e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=11e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=11e-6
m7 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=99e-6
m8 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=174e-6
m9 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=68e-6
m10 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=5e-6 W=183e-6
m11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
m13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=153e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=18e-6
m15 outFirstStage outInputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=521e-6
m16 out outInputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=564e-6
m17 FirstStageYout1 outInputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=521e-6
m18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=33e-6
m19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=33e-6
m20 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=224e-6
Capacitor1 outFirstStage out 13.9001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_78_3

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 5.08301 mW
** Area: 12930 (mu_m)^2
** Transit frequency: 2.69201 MHz
** Transit frequency with error factor: 2.69162 MHz
** Slew rate: 4.98555 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 3.22001 V
** VoutMin: 0.550001 V
** VcmMax: 4.66001 V
** VcmMin: 1.62001 V


** Expected Currents: 
** NormalTransistorNmos: 3.72281e+07 muA
** NormalTransistorPmos: -7.00259e+07 muA
** NormalTransistorPmos: -1.11686e+08 muA
** NormalTransistorPmos: -7.00259e+07 muA
** NormalTransistorPmos: -1.11686e+08 muA
** DiodeTransistorNmos: 7.00251e+07 muA
** DiodeTransistorNmos: 7.00241e+07 muA
** NormalTransistorNmos: 7.00251e+07 muA
** NormalTransistorNmos: 7.00241e+07 muA
** NormalTransistorNmos: 8.33251e+07 muA
** DiodeTransistorNmos: 8.33261e+07 muA
** NormalTransistorNmos: 4.16621e+07 muA
** NormalTransistorNmos: 4.16621e+07 muA
** NormalTransistorNmos: 7.45974e+08 muA
** NormalTransistorPmos: -7.45973e+08 muA
** NormalTransistorPmos: -7.45974e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.72289e+07 muA
** DiodeTransistorPmos: -3.72289e+07 muA


** Expected Voltages: 
** ibias: 1.26401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.959001  V
** outInputVoltageBiasXXpXX1: 2.37201  V
** outSourceVoltageBiasXXnXX1: 0.633001  V
** outSourceVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.554001  V
** out1: 1.16401  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.74301  V
** innerStageBias: 3.40501  V
** inner: 0.629001  V


.END