.suckt  one_stage_fully_differential_op_amp16 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m5 outFeedback outFeedback sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX1 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m7 FeedbackStageYinnerStageBias1 ibias sourceNmos sourceNmos nmos
m8 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX1 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m9 FeedbackStageYinnerStageBias2 ibias sourceNmos sourceNmos nmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m14 out1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m15 FirstStageYinnerTransistorStack1Load1 outFeedback sourcePmos sourcePmos pmos
m16 out2 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m17 FirstStageYinnerTransistorStack2Load1 outFeedback sourcePmos sourcePmos pmos
m18 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m19 out1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m20 out2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out1 sourceNmos 
c2 out2 sourceNmos 
m21 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m22 ibias ibias sourceNmos sourceNmos nmos
m23 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m24 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end one_stage_fully_differential_op_amp16

