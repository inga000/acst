.suckt  symmetrical_op_amp85 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage out2FirstStage out1FirstStage out1FirstStage nmos
m2 out1FirstStage out1FirstStage sourceNmos sourceNmos nmos
m3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage nmos
m4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m5 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m6 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m7 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c1 out sourceNmos 
m8 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m9 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m10 out innerComplementarySecondStage sourcePmos sourcePmos pmos
m11 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos
m12 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m13 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m14 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp85

