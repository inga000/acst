** Name: two_stage_single_output_op_amp_19_2

.MACRO two_stage_single_output_op_amp_19_2 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=73e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=32e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=32e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=214e-6
mMainBias8 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=209e-6
mSecondStage1Transconductor9 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=76e-6
mSimpleFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=7e-6
mSimpleFirstStageStageBias11 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=76e-6
mSimpleFirstStageTransconductor12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=14e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=4e-6 W=167e-6
mSecondStage1StageBias14 out ibias sourcePmos sourcePmos pmos4 L=6e-6 W=322e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=14e-6
mMainBias16 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=89e-6
mMainBias17 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=82e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_19_2

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 1.40201 mW
** Area: 7014 (mu_m)^2
** Transit frequency: 2.74501 MHz
** Transit frequency with error factor: 2.74074 MHz
** Slew rate: 4.16286 V/mu_s
** Phase margin: 63.5984°
** CMRR: 100 dB
** negPSRR: 100 dB
** posPSRR: 115 dB
** VoutMax: 4.68001 V
** VoutMin: 0.330001 V
** VcmMax: 3.06001 V
** VcmMin: 0.190001 V


** Expected Currents: 
** NormalTransistorNmos: 7.98801e+07 muA
** NormalTransistorPmos: -2.82809e+07 muA
** NormalTransistorPmos: -2.58479e+07 muA
** DiodeTransistorNmos: 1.20631e+07 muA
** NormalTransistorNmos: 1.20631e+07 muA
** NormalTransistorNmos: 1.20631e+07 muA
** NormalTransistorPmos: -2.41289e+07 muA
** NormalTransistorPmos: -2.41299e+07 muA
** NormalTransistorPmos: -1.20639e+07 muA
** NormalTransistorPmos: -1.20639e+07 muA
** NormalTransistorNmos: 1.0232e+08 muA
** NormalTransistorNmos: 1.02319e+08 muA
** NormalTransistorPmos: -1.02319e+08 muA
** DiodeTransistorNmos: 2.82801e+07 muA
** DiodeTransistorNmos: 2.58471e+07 muA
** DiodeTransistorPmos: -7.98809e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.11101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.556001  V
** outVoltageBiasXXnXX1: 0.756001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.42901  V
** innerTransistorStack2Load1: 0.150001  V
** out1: 0.555001  V
** sourceTransconductance: 3.37301  V
** innerTransconductance: 0.172001  V


.END