.suckt  two_stage_single_output_op_amp_1_8 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad3 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias7 out outInputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
mSecondStage1StageBias8 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mSecondStage1Transconductor9 out outFirstStage sourcePmos sourcePmos pmos
mMainBias10 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mMainBias11 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias12 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_1_8

