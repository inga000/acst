** Name: two_stage_single_output_op_amp_8_8

.MACRO two_stage_single_output_op_amp_8_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=19e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=107e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=6e-6 W=106e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=600e-6
mSecondStage1StageBias8 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=7e-6 W=93e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=10e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=19e-6
mMainBias11 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=35e-6
mSecondStage1Transconductor12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=411e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=107e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_8_8

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 2.18801 mW
** Area: 6581 (mu_m)^2
** Transit frequency: 5.32601 MHz
** Transit frequency with error factor: 5.3179 MHz
** Slew rate: 6.04009 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** negPSRR: 157 dB
** posPSRR: 97 dB
** VoutMax: 4.79001 V
** VoutMin: 0.720001 V
** VcmMax: 4.63001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorNmos: 9.88701e+06 muA
** NormalTransistorPmos: -4.40659e+07 muA
** DiodeTransistorPmos: -2.75779e+07 muA
** NormalTransistorPmos: -2.75779e+07 muA
** NormalTransistorNmos: 5.51541e+07 muA
** NormalTransistorNmos: 2.75771e+07 muA
** NormalTransistorNmos: 2.75771e+07 muA
** NormalTransistorNmos: 3.18499e+08 muA
** NormalTransistorNmos: 3.18498e+08 muA
** NormalTransistorPmos: -3.18498e+08 muA
** DiodeTransistorNmos: 4.40651e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.88799e+06 muA


** Expected Voltages: 
** ibias: 0.598001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.12801  V
** out: 2.5  V
** outFirstStage: 4.22701  V
** outVoltageBiasXXpXX0: 3.68901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.22701  V
** sourceTransconductance: 1.91401  V
** innerStageBias: 0.193001  V


.END