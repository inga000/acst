.suckt  two_stage_fully_differential_op_amp_13_7 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m2 outFeedback outFeedback sourcePmos sourcePmos pmos
m3 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m4 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m5 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m6 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m7 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m8 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m9 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m10 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m12 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m13 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m14 out1 ibias sourceNmos sourceNmos nmos
m15 out1 out1FirstStage sourcePmos sourcePmos pmos
m16 out2 ibias sourceNmos sourceNmos nmos
m17 out2 out2FirstStage sourcePmos sourcePmos pmos
m18 ibias ibias sourceNmos sourceNmos nmos
.end two_stage_fully_differential_op_amp_13_7

