** Name: two_stage_single_output_op_amp_58_12

.MACRO two_stage_single_output_op_amp_58_12 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=18e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=18e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=178e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=75e-6
m5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=24e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=564e-6
m7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
m8 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=63e-6
m9 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=178e-6
m10 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=156e-6
m11 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=156e-6
m12 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=156e-6
m13 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=292e-6
m14 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=292e-6
m15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
m16 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=174e-6
m17 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=598e-6
m18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=63e-6
m19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=359e-6
m20 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=453e-6
m21 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=453e-6
m22 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=564e-6
m23 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=599e-6
m24 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=24e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 13.6001e-12
.EOM two_stage_single_output_op_amp_58_12

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 12.4281 mW
** Area: 14975 (mu_m)^2
** Transit frequency: 9.35201 MHz
** Transit frequency with error factor: 9.3385 MHz
** Slew rate: 12.2242 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 1.30001 V
** VcmMax: 3.04001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.52301e+08 muA
** NormalTransistorPmos: -1.50718e+08 muA
** NormalTransistorPmos: -7.26169e+07 muA
** NormalTransistorNmos: 1.66817e+08 muA
** NormalTransistorNmos: 2.85973e+08 muA
** NormalTransistorNmos: 1.66815e+08 muA
** NormalTransistorNmos: 2.85969e+08 muA
** DiodeTransistorPmos: -1.66814e+08 muA
** NormalTransistorPmos: -1.66814e+08 muA
** NormalTransistorPmos: -2.38308e+08 muA
** DiodeTransistorPmos: -2.38307e+08 muA
** NormalTransistorPmos: -1.19154e+08 muA
** NormalTransistorPmos: -1.19154e+08 muA
** NormalTransistorNmos: 1.51794e+09 muA
** DiodeTransistorNmos: 1.51794e+09 muA
** NormalTransistorPmos: -1.51793e+09 muA
** NormalTransistorPmos: -1.51793e+09 muA
** DiodeTransistorNmos: 1.50719e+08 muA
** NormalTransistorNmos: 1.50719e+08 muA
** DiodeTransistorNmos: 7.26161e+07 muA
** DiodeTransistorNmos: 7.26151e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.523e+08 muA


** Expected Voltages: 
** ibias: 3.34001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.27001  V
** out: 2.5  V
** outFirstStage: 4.06101  V
** outInputVoltageBiasXXnXX1: 1.70401  V
** outSourceVoltageBiasXXnXX1: 0.852001  V
** outSourceVoltageBiasXXnXX2: 0.557001  V
** outSourceVoltageBiasXXpXX1: 4.17101  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.05001  V
** sourceGCC1: 0.706001  V
** sourceGCC2: 0.706001  V
** sourceTransconductance: 3.36001  V
** innerTransconductance: 4.625  V
** inner: 0.852001  V
** inner: 4.16801  V


.END