** Name: two_stage_single_output_op_amp_52_5

.MACRO two_stage_single_output_op_amp_52_5 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
m2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=293e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=26e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=73e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=574e-6
m7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=320e-6
m8 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=239e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=516e-6
m10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=32e-6
m11 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=114e-6
m12 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=293e-6
m13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=301e-6
m14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=301e-6
m15 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=145e-6
m16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=352e-6
m17 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=574e-6
m18 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=12e-6
m19 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=12e-6
m20 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=235e-6
m21 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=235e-6
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=73e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 7e-12
.EOM two_stage_single_output_op_amp_52_5

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 10.2521 mW
** Area: 14995 (mu_m)^2
** Transit frequency: 21.5541 MHz
** Transit frequency with error factor: 21.5537 MHz
** Slew rate: 15.9095 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 3.36001 V
** VoutMin: 0.150001 V
** VcmMax: 5.19001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorNmos: 1.25376e+08 muA
** NormalTransistorNmos: 2.63988e+08 muA
** NormalTransistorPmos: -2.85583e+08 muA
** NormalTransistorPmos: -1.11626e+08 muA
** NormalTransistorPmos: -1.91361e+08 muA
** NormalTransistorPmos: -1.11625e+08 muA
** NormalTransistorPmos: -1.9136e+08 muA
** DiodeTransistorNmos: 1.11627e+08 muA
** NormalTransistorNmos: 1.11626e+08 muA
** NormalTransistorNmos: 1.11627e+08 muA
** NormalTransistorNmos: 1.5947e+08 muA
** NormalTransistorNmos: 7.97341e+07 muA
** NormalTransistorNmos: 7.97341e+07 muA
** NormalTransistorNmos: 9.82788e+08 muA
** NormalTransistorPmos: -9.82787e+08 muA
** DiodeTransistorPmos: -9.82788e+08 muA
** DiodeTransistorNmos: 2.85584e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.25375e+08 muA
** NormalTransistorPmos: -1.25376e+08 muA
** DiodeTransistorPmos: -2.63987e+08 muA
** DiodeTransistorPmos: -2.63988e+08 muA


** Expected Voltages: 
** ibias: 0.567001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.957001  V
** inputVoltageBiasXXpXX2: 2.90801  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.79601  V
** outSourceVoltageBiasXXpXX1: 3.89801  V
** outSourceVoltageBiasXXpXX2: 4.22201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.19001  V
** sourceGCC2: 4.19001  V
** sourceTransconductance: 1.92701  V
** inner: 3.89501  V


.END