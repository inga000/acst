.suckt  symmetrical_op_amp33 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_MainBias_1 inOutputStageBiasComplementarySecondStage outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_3 outFirstStage outFirstStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Load_4 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_StageBias_5 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m_Symmetrical_FirstStage_StageBias_6 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Transconductor_7 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_Symmetrical_FirstStage_Transconductor_8 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_Transconductor_9 out outFirstStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_StageBias_10 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m_Symmetrical_SecondStage1_StageBias_11 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_12 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_13 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_14 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_15 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_16 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_MainBias_17 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp33

