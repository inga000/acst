** Name: two_stage_single_output_op_amp_190_9

.MACRO two_stage_single_output_op_amp_190_9 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=352e-6
m2 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=1e-6 W=13e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=27e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=248e-6
m5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=25e-6
m6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=61e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=10e-6
m8 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=30e-6
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=6e-6
m10 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=248e-6
m11 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=25e-6
m12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=6e-6
m13 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=27e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=352e-6
m15 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
m16 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=385e-6
m17 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=140e-6
m18 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=204e-6
m19 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=25e-6
m20 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=126e-6
m21 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=126e-6
m22 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=385e-6
Capacitor1 outFirstStage out 4.5e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_190_9

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 4.91001 mW
** Area: 14332 (mu_m)^2
** Transit frequency: 2.54601 MHz
** Transit frequency with error factor: 2.54379 MHz
** Slew rate: 3.50006 V/mu_s
** Phase margin: 62.4525°
** CMRR: 117 dB
** VoutMax: 4.25 V
** VoutMin: 0.700001 V
** VcmMax: 4.57001 V
** VcmMin: 1.5 V


** Expected Currents: 
** NormalTransistorPmos: -2.07135e+08 muA
** NormalTransistorPmos: -2.50119e+07 muA
** NormalTransistorNmos: 1.19946e+08 muA
** NormalTransistorNmos: 1.19947e+08 muA
** DiodeTransistorNmos: 1.19946e+08 muA
** NormalTransistorPmos: -1.28047e+08 muA
** NormalTransistorPmos: -1.28048e+08 muA
** NormalTransistorPmos: -1.28048e+08 muA
** NormalTransistorPmos: -1.28048e+08 muA
** NormalTransistorNmos: 1.62051e+07 muA
** DiodeTransistorNmos: 1.62041e+07 muA
** NormalTransistorNmos: 8.10201e+06 muA
** NormalTransistorNmos: 8.10201e+06 muA
** NormalTransistorNmos: 4.73825e+08 muA
** DiodeTransistorNmos: 4.73824e+08 muA
** NormalTransistorPmos: -4.73824e+08 muA
** DiodeTransistorNmos: 2.07136e+08 muA
** NormalTransistorNmos: 2.07137e+08 muA
** DiodeTransistorNmos: 2.50111e+07 muA
** NormalTransistorNmos: 2.50101e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.12601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.28401  V
** outInputVoltageBiasXXnXX2: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.642001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.90501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 3.99401  V
** innerTransistorStack2Load1: 1.15501  V
** innerTransistorStack2Load2: 3.99401  V
** out1: 2.09501  V
** sourceTransconductance: 1.87601  V
** inner: 0.643001  V
** inner: 0.554001  V


.END