** Name: two_stage_single_output_op_amp_53_8

.MACRO two_stage_single_output_op_amp_53_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=13e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=21e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=197e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=52e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=52e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=441e-6
mSecondStage1StageBias12 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=8e-6 W=576e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=84e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=50e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=50e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=276e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=84e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=126e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=414e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.10001e-12
.EOM two_stage_single_output_op_amp_53_8

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 7.97001 mW
** Area: 8180 (mu_m)^2
** Transit frequency: 5.35301 MHz
** Transit frequency with error factor: 5.35335 MHz
** Slew rate: 6.59022 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.550001 V
** VcmMax: 5.17001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorPmos: -1.26253e+08 muA
** NormalTransistorPmos: -4.1218e+08 muA
** NormalTransistorPmos: -3.37959e+07 muA
** NormalTransistorPmos: -5.06929e+07 muA
** NormalTransistorPmos: -3.37959e+07 muA
** NormalTransistorPmos: -5.06929e+07 muA
** DiodeTransistorNmos: 3.37951e+07 muA
** DiodeTransistorNmos: 3.37941e+07 muA
** NormalTransistorNmos: 3.37951e+07 muA
** NormalTransistorNmos: 3.37941e+07 muA
** NormalTransistorNmos: 3.37951e+07 muA
** NormalTransistorNmos: 1.68981e+07 muA
** NormalTransistorNmos: 1.68981e+07 muA
** NormalTransistorNmos: 9.34113e+08 muA
** NormalTransistorNmos: 9.34112e+08 muA
** NormalTransistorPmos: -9.34112e+08 muA
** DiodeTransistorNmos: 1.26254e+08 muA
** DiodeTransistorNmos: 4.12181e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.15501  V
** outVoltageBiasXXnXX2: 0.563001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.574001  V
** innerTransistorStack2Load2: 0.573001  V
** out1: 1.15401  V
** sourceGCC1: 4.11201  V
** sourceGCC2: 4.11201  V
** sourceTransconductance: 1.89901  V
** innerStageBias: 0.358001  V


.END