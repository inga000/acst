** Name: two_stage_single_output_op_amp_1_3

.MACRO two_stage_single_output_op_amp_1_3 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=184e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=11e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=5e-6
m5 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=363e-6
m6 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=184e-6
m7 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=12e-6
m8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=19e-6
m9 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=127e-6
m10 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=252e-6
m11 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=5e-6 W=469e-6
m12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=19e-6
m13 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_1_3

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 1.93701 mW
** Area: 6799 (mu_m)^2
** Transit frequency: 5.67501 MHz
** Transit frequency with error factor: 5.64444 MHz
** Slew rate: 9.38409 V/mu_s
** Phase margin: 67.0361°
** CMRR: 88 dB
** negPSRR: 89 dB
** posPSRR: 208 dB
** VoutMax: 4.31001 V
** VoutMin: 0.150001 V
** VcmMax: 3.40001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 1.01161e+07 muA
** NormalTransistorPmos: -8.31699e+06 muA
** DiodeTransistorNmos: 5.86851e+07 muA
** NormalTransistorNmos: 5.86851e+07 muA
** NormalTransistorPmos: -1.1737e+08 muA
** NormalTransistorPmos: -5.86859e+07 muA
** NormalTransistorPmos: -5.86859e+07 muA
** NormalTransistorNmos: 2.31554e+08 muA
** NormalTransistorPmos: -2.31553e+08 muA
** NormalTransistorPmos: -2.31554e+08 muA
** DiodeTransistorNmos: 8.31601e+06 muA
** DiodeTransistorPmos: -1.01169e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.11601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.719001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceTransconductance: 3.78101  V
** innerStageBias: 4.62001  V


.END