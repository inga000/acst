.suckt  two_stage_single_output_op_amp_152_5 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mMainBias2 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad5 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad9 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSimpleFirstStageTransconductor12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1Transconductor14 out outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias15 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mSecondStage1StageBias16 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mMainBias17 ibias ibias sourceNmos sourceNmos nmos
mMainBias18 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mMainBias20 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
mMainBias21 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_152_5

