.suckt  two_stage_single_output_op_amp_189_4 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_2 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_3 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_4 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m_SingleOutput_FirstStage_Load_5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_6 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m_SingleOutput_FirstStage_Load_7 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_8 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m_SingleOutput_FirstStage_Load_9 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_StageBias_10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_SingleOutput_FirstStage_StageBias_11 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Transconductor_12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_SingleOutput_FirstStage_Transconductor_13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_Transconductor_14 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_SingleOutput_SecondStage1_Transconductor_15 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_16 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m_SingleOutput_SecondStage1_StageBias_17 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_SecondStage1_StageBias_18 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_19 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_20 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_SingleOutput_MainBias_21 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_189_4

