.suckt  two_stage_single_output_op_amp_136_10 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias2 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mMainBias3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mSimpleFirstStageLoad4 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad6 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias15 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSecondStage1Transconductor16 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
mMainBias18 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias19 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias20 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mMainBias21 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_136_10

