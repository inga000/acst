** Name: two_stage_single_output_op_amp_47_9

.MACRO two_stage_single_output_op_amp_47_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=10e-6 W=13e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=15e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=287e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=11e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=8e-6 W=146e-6
mMainBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=10e-6 W=39e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=63e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=63e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=287e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=10e-6 W=39e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=140e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=35e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=35e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=14e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=14e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=8e-6 W=519e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=108e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=598e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=140e-6
mMainBias23 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=415e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_47_9

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 3.47701 mW
** Area: 14974 (mu_m)^2
** Transit frequency: 2.70601 MHz
** Transit frequency with error factor: 2.70562 MHz
** Slew rate: 5.51797 V/mu_s
** Phase margin: 71.0468°
** CMRR: 130 dB
** VoutMax: 4.68001 V
** VoutMin: 0.700001 V
** VcmMax: 3.80001 V
** VcmMin: -0.279999 V


** Expected Currents: 
** NormalTransistorNmos: 6.84801e+06 muA
** NormalTransistorPmos: -2.85709e+07 muA
** NormalTransistorPmos: -7.38399e+06 muA
** NormalTransistorNmos: 2.51031e+07 muA
** NormalTransistorNmos: 4.30351e+07 muA
** NormalTransistorNmos: 2.50991e+07 muA
** NormalTransistorNmos: 4.30291e+07 muA
** NormalTransistorPmos: -2.51019e+07 muA
** NormalTransistorPmos: -2.51009e+07 muA
** NormalTransistorPmos: -2.50999e+07 muA
** NormalTransistorPmos: -2.51009e+07 muA
** NormalTransistorPmos: -3.58619e+07 muA
** NormalTransistorPmos: -1.79309e+07 muA
** NormalTransistorPmos: -1.79309e+07 muA
** NormalTransistorNmos: 5.46629e+08 muA
** DiodeTransistorNmos: 5.46629e+08 muA
** NormalTransistorPmos: -5.46628e+08 muA
** DiodeTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** DiodeTransistorNmos: 7.38301e+06 muA
** DiodeTransistorNmos: 7.38401e+06 muA
** DiodeTransistorPmos: -6.84899e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.35101  V
** inputVoltageBiasXXpXX1: 3.81401  V
** out: 2.5  V
** outFirstStage: 4.11501  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.688001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.23501  V
** innerTransistorStack1Load2: 4.57801  V
** innerTransistorStack2Load2: 4.57801  V
** sourceGCC1: 0.669001  V
** sourceGCC2: 0.669001  V
** sourceTransconductance: 3.52601  V
** inner: 0.555001  V


.END