** Name: symmetrical_op_amp188

.MACRO symmetrical_op_amp188 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=10e-6
mSecondStage1StageBias2 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=8e-6 W=108e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias4 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mSymmetricalFirstStageStageBias5 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=48e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=21e-6
mSymmetricalFirstStageTransconductor7 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=42e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias8 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=8e-6 W=108e-6
mSecondStage1StageBias9 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos4 L=2e-6 W=42e-6
mSymmetricalFirstStageTransconductor10 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=42e-6
mMainBias11 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=38e-6
mSymmetricalFirstStageLoad12 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=10e-6
mSymmetricalFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=10e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=30e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=30e-6
mSymmetricalFirstStageLoad16 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=79e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=241e-6
mSecondStage1Transconductor18 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=241e-6
mSymmetricalFirstStageLoad19 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=79e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp188

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 0.824001 mW
** Area: 4238 (mu_m)^2
** Transit frequency: 5.07701 MHz
** Transit frequency with error factor: 5.07703 MHz
** Slew rate: 4.85868 V/mu_s
** Phase margin: 77.9223°
** CMRR: 144 dB
** negPSRR: 130 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 0.780001 V
** VcmMax: 4.81001 V
** VcmMin: 1.35001 V


** Expected Currents: 
** NormalTransistorNmos: 2.53531e+07 muA
** NormalTransistorPmos: -1.6e+07 muA
** NormalTransistorPmos: -1.60009e+07 muA
** NormalTransistorPmos: -1.6e+07 muA
** NormalTransistorPmos: -1.60009e+07 muA
** NormalTransistorNmos: 3.19971e+07 muA
** NormalTransistorNmos: 3.19961e+07 muA
** NormalTransistorNmos: 1.59991e+07 muA
** NormalTransistorNmos: 1.59991e+07 muA
** NormalTransistorNmos: 4.87361e+07 muA
** DiodeTransistorNmos: 4.87351e+07 muA
** NormalTransistorPmos: -4.87369e+07 muA
** NormalTransistorPmos: -4.87359e+07 muA
** NormalTransistorNmos: 4.87361e+07 muA
** NormalTransistorPmos: -4.87369e+07 muA
** NormalTransistorPmos: -4.87359e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.53539e+07 muA


** Expected Voltages: 
** ibias: 1.15101  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** inStageBiasComplementarySecondStage: 0.611001  V
** innerComplementarySecondStage: 1.18101  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.513001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END