** Name: two_stage_single_output_op_amp_19_5

.MACRO two_stage_single_output_op_amp_19_5 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=173e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=51e-6
m3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
m4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=101e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=133e-6
m7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=173e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=323e-6
m10 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=27e-6
m11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=428e-6
m12 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=530e-6
m13 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=93e-6
m14 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=47e-6
m15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=101e-6
m16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=133e-6
m17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=530e-6
m18 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=55e-6
m19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_19_5

** Expected Performance Values: 
** Gain: 106 dB
** Power consumption: 6.42401 mW
** Area: 14085 (mu_m)^2
** Transit frequency: 16.3121 MHz
** Transit frequency with error factor: 16.2977 MHz
** Slew rate: 20.4529 V/mu_s
** Phase margin: 65.3172°
** CMRR: 104 dB
** negPSRR: 106 dB
** posPSRR: 228 dB
** VoutMax: 3 V
** VoutMin: 0.150001 V
** VcmMax: 3.10001 V
** VcmMin: 0.370001 V


** Expected Currents: 
** NormalTransistorNmos: 4.71236e+08 muA
** NormalTransistorPmos: -5.57629e+07 muA
** NormalTransistorPmos: -2.73469e+07 muA
** DiodeTransistorNmos: 4.71451e+07 muA
** NormalTransistorNmos: 4.71451e+07 muA
** NormalTransistorNmos: 4.71451e+07 muA
** NormalTransistorPmos: -9.42909e+07 muA
** NormalTransistorPmos: -9.42899e+07 muA
** NormalTransistorPmos: -4.71459e+07 muA
** NormalTransistorPmos: -4.71459e+07 muA
** NormalTransistorNmos: 6.16168e+08 muA
** NormalTransistorPmos: -6.16167e+08 muA
** DiodeTransistorPmos: -6.16168e+08 muA
** DiodeTransistorNmos: 5.57621e+07 muA
** DiodeTransistorNmos: 2.73461e+07 muA
** DiodeTransistorPmos: -4.71235e+08 muA
** NormalTransistorPmos: -4.71235e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.43601  V
** outSourceVoltageBiasXXpXX1: 3.71701  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.602001  V
** outVoltageBiasXXnXX1: 0.934001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerStageBias: 4.29601  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.26301  V
** inner: 3.71901  V


.END