.suckt  symmetrical_op_amp39 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_FirstStage_Load_1 outFirstStage outFirstStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Load_2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_StageBias_3 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m_Symmetrical_FirstStage_StageBias_4 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Transconductor_5 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_Symmetrical_FirstStage_Transconductor_6 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage2_Transconductor_7 out outFirstStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage2_StageBias_8 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos
m_Symmetrical_SecondStage2_StageBias_9 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_10 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_11 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_12 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_Symmetrical_MainBias_13 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end symmetrical_op_amp39

