** Name: two_stage_single_output_op_amp_143_8

.MACRO two_stage_single_output_op_amp_143_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=19e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=42e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=381e-6
mSecondStage1StageBias9 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=368e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=11e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=42e-6
mSimpleFirstStageLoad12 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=181e-6
mMainBias13 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=220e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=212e-6
mSimpleFirstStageLoad15 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=181e-6
mMainBias16 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=548e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.2001e-12
.EOM two_stage_single_output_op_amp_143_8

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 14.1971 mW
** Area: 2855 (mu_m)^2
** Transit frequency: 6.92501 MHz
** Transit frequency with error factor: 6.91241 MHz
** Slew rate: 6.527 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 0.630001 V
** VcmMax: 5.22001 V
** VcmMin: 0.810001 V


** Expected Currents: 
** NormalTransistorPmos: -3.24451e+08 muA
** NormalTransistorPmos: -1.29311e+08 muA
** NormalTransistorNmos: 6.65271e+07 muA
** NormalTransistorNmos: 6.65281e+07 muA
** DiodeTransistorNmos: 6.65271e+07 muA
** NormalTransistorPmos: -1.06525e+08 muA
** NormalTransistorPmos: -1.06525e+08 muA
** NormalTransistorNmos: 7.99951e+07 muA
** NormalTransistorNmos: 3.99981e+07 muA
** NormalTransistorNmos: 3.99981e+07 muA
** NormalTransistorNmos: 2.15253e+09 muA
** NormalTransistorNmos: 2.15253e+09 muA
** NormalTransistorPmos: -2.15252e+09 muA
** DiodeTransistorNmos: 3.24452e+08 muA
** DiodeTransistorNmos: 1.29312e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.664001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 1.03701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** out1: 2.21801  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.259001  V


.END