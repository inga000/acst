** Name: two_stage_single_output_op_amp_71_4

.MACRO two_stage_single_output_op_amp_71_4 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=34e-6
mSecondStage1StageBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=418e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=37e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=24e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=24e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=19e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=270e-6
mSecondStage1Transconductor11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=178e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=34e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=122e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=11e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=11e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=101e-6
mSecondStage1StageBias17 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=596e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=122e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=64e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=130e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_71_4

** Expected Performance Values: 
** Gain: 148 dB
** Power consumption: 4.13601 mW
** Area: 6900 (mu_m)^2
** Transit frequency: 4.38701 MHz
** Transit frequency with error factor: 4.3841 MHz
** Slew rate: 3.64262 V/mu_s
** Phase margin: 60.7336°
** CMRR: 108 dB
** VoutMax: 3.52001 V
** VoutMin: 0.330001 V
** VcmMax: 4.75 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorPmos: -1.62037e+08 muA
** NormalTransistorPmos: -3.31491e+08 muA
** NormalTransistorPmos: -1.65159e+07 muA
** NormalTransistorPmos: -2.80489e+07 muA
** NormalTransistorPmos: -1.65159e+07 muA
** NormalTransistorPmos: -2.80489e+07 muA
** DiodeTransistorNmos: 1.65151e+07 muA
** NormalTransistorNmos: 1.65151e+07 muA
** NormalTransistorNmos: 2.30631e+07 muA
** NormalTransistorNmos: 2.30621e+07 muA
** NormalTransistorNmos: 1.15321e+07 muA
** NormalTransistorNmos: 1.15321e+07 muA
** NormalTransistorNmos: 2.57544e+08 muA
** NormalTransistorNmos: 2.57543e+08 muA
** NormalTransistorPmos: -2.57543e+08 muA
** NormalTransistorPmos: -2.57542e+08 muA
** DiodeTransistorNmos: 1.62038e+08 muA
** DiodeTransistorNmos: 3.31492e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.00701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.78501  V
** outVoltageBiasXXnXX1: 0.967001  V
** outVoltageBiasXXnXX2: 0.598001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.393001  V
** out1: 0.556001  V
** sourceGCC1: 3.72101  V
** sourceGCC2: 3.72101  V
** sourceTransconductance: 1.91001  V
** innerStageBias: 3.83901  V
** innerTransconductance: 0.377001  V


.END