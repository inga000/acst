** Name: two_stage_single_output_op_amp_11_8

.MACRO two_stage_single_output_op_amp_11_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=7e-6 W=61e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=7e-6 W=47e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=52e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=14e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=14e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=345e-6
mMainBias9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=32e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=283e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=14e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=7e-6 W=47e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=203e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=7e-6 W=61e-6
mMainBias15 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=29e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_11_8

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 4.11301 mW
** Area: 4855 (mu_m)^2
** Transit frequency: 2.84001 MHz
** Transit frequency with error factor: 2.83696 MHz
** Slew rate: 6.07411 V/mu_s
** Phase margin: 70.4739°
** CMRR: 97 dB
** negPSRR: 93 dB
** posPSRR: 87 dB
** VoutMax: 4.25 V
** VoutMin: 0.560001 V
** VcmMax: 3.64001 V
** VcmMin: 1.01001 V


** Expected Currents: 
** NormalTransistorNmos: 6.33671e+07 muA
** NormalTransistorPmos: -3.46719e+07 muA
** DiodeTransistorPmos: -1.37339e+07 muA
** DiodeTransistorPmos: -1.37349e+07 muA
** NormalTransistorPmos: -1.37339e+07 muA
** NormalTransistorPmos: -1.37349e+07 muA
** NormalTransistorNmos: 2.74671e+07 muA
** NormalTransistorNmos: 1.37331e+07 muA
** NormalTransistorNmos: 1.37331e+07 muA
** NormalTransistorNmos: 6.87047e+08 muA
** NormalTransistorNmos: 6.87046e+08 muA
** NormalTransistorPmos: -6.87046e+08 muA
** DiodeTransistorNmos: 3.46711e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.33679e+07 muA


** Expected Voltages: 
** ibias: 0.670001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.85501  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 0.962001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.23801  V
** innerTransistorStack1Load1: 4.09801  V
** innerTransistorStack2Load1: 4.09801  V
** sourceTransconductance: 1.75301  V
** innerStageBias: 0.265001  V


.END