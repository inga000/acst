.suckt  symmetrical_op_amp16 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m3 outFirstStage outFirstStage sourcePmos sourcePmos pmos
m4 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m6 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m7 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m8 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m9 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
m10 out outFirstStage sourcePmos sourcePmos pmos
m11 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
m12 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m13 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m14 ibias ibias sourceNmos sourceNmos nmos
m15 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end symmetrical_op_amp16

