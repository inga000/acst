** Name: one_stage_single_output_op_amp101

.MACRO one_stage_single_output_op_amp101 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
m2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=19e-6
m4 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
m5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=7e-6
m6 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=40e-6
m7 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m8 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m9 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=192e-6
m10 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
m11 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=597e-6
m12 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=79e-6
m13 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=192e-6
m14 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=340e-6
m15 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=340e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp101

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 0.955001 mW
** Area: 6949 (mu_m)^2
** Transit frequency: 5.40001 MHz
** Transit frequency with error factor: 5.40013 MHz
** Slew rate: 8.0168 V/mu_s
** Phase margin: 63.0254°
** CMRR: 145 dB
** VoutMax: 3.17001 V
** VoutMin: 0.850001 V
** VcmMax: 3 V
** VcmMin: 0.690001 V


** Expected Currents: 
** NormalTransistorNmos: 8.27401e+06 muA
** NormalTransistorPmos: -1.00569e+07 muA
** NormalTransistorPmos: -7.62979e+07 muA
** NormalTransistorPmos: -7.62989e+07 muA
** NormalTransistorNmos: 7.62971e+07 muA
** NormalTransistorNmos: 7.62981e+07 muA
** DiodeTransistorNmos: 7.62971e+07 muA
** NormalTransistorPmos: -1.60869e+08 muA
** NormalTransistorPmos: -1.60868e+08 muA
** NormalTransistorPmos: -7.62979e+07 muA
** NormalTransistorPmos: -7.62979e+07 muA
** DiodeTransistorNmos: 1.00561e+07 muA
** DiodeTransistorPmos: -8.27499e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.15401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX2: 3.96101  V
** outVoltageBiasXXnXX0: 0.603001  V
** outVoltageBiasXXpXX1: 2.04501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.28701  V
** innerSourceLoad2: 0.704001  V
** innerStageBias: 3.89101  V
** out1: 1.25901  V
** sourceGCC1: 3.00501  V
** sourceGCC2: 3.00501  V


.END