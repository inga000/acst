.suckt  symmetrical_op_amp15 ibias in1 in2 out sourceNmos sourcePmos
m1 outFirstStage outFirstStage sourcePmos sourcePmos pmos
m2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m3 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m4 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m5 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m6 out innerComplementarySecondStage sourceNmos sourceNmos nmos
m7 out outFirstStage sourcePmos sourcePmos pmos
m8 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
m9 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m10 ibias ibias sourceNmos sourceNmos nmos
.end symmetrical_op_amp15

