.suckt  two_stage_fully_differential_op_amp_5_8 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m3 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m4 outFeedback outFeedback sourceNmos sourceNmos nmos
m5 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m7 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m8 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m9 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m10 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m11 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m12 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m13 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m14 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m15 out1FirstStage ibias sourcePmos sourcePmos pmos
m16 out2FirstStage ibias sourcePmos sourcePmos pmos
m17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m20 out1 outVoltageBiasXXnXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias nmos
m21 SecondStage1YinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m22 out1 out1FirstStage sourcePmos sourcePmos pmos
m23 out2 outVoltageBiasXXnXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias nmos
m24 SecondStage2YinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m25 out2 out2FirstStage sourcePmos sourcePmos pmos
m26 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m27 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m28 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_5_8

