** Name: two_stage_single_output_op_amp_10_7

.MACRO two_stage_single_output_op_amp_10_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=15e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=10e-6 W=24e-6
mSimpleFirstStageTransconductor4 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=20e-6
mSimpleFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
mMainBias6 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mSecondStage1StageBias7 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=233e-6
mSimpleFirstStageTransconductor8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=20e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=15e-6
mSecondStage1Transconductor10 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=75e-6
mSimpleFirstStageLoad11 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=10e-6 W=192e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_10_7

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 2.55301 mW
** Area: 3552 (mu_m)^2
** Transit frequency: 3.51901 MHz
** Transit frequency with error factor: 3.51606 MHz
** Slew rate: 3.94978 V/mu_s
** Phase margin: 62.4525°
** CMRR: 97 dB
** negPSRR: 137 dB
** posPSRR: 95 dB
** VoutMax: 4.42001 V
** VoutMin: 0.260001 V
** VcmMax: 4.10001 V
** VcmMin: 0.850001 V


** Expected Currents: 
** NormalTransistorNmos: 2.40181e+07 muA
** DiodeTransistorPmos: -9.00799e+06 muA
** NormalTransistorPmos: -9.00799e+06 muA
** NormalTransistorPmos: -9.00799e+06 muA
** NormalTransistorNmos: 1.80131e+07 muA
** NormalTransistorNmos: 9.00701e+06 muA
** NormalTransistorNmos: 9.00701e+06 muA
** NormalTransistorNmos: 4.5856e+08 muA
** NormalTransistorPmos: -4.58559e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.40189e+07 muA


** Expected Voltages: 
** ibias: 0.670001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.85401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.41201  V
** out1: 3.85401  V
** sourceTransconductance: 1.91601  V


.END