** Name: symmetrical_op_amp37

.MACRO symmetrical_op_amp37 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=9e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias4 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=111e-6
mMainBias6 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
mMainBias9 inOutputStageBiasComplementarySecondStage outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=51e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=95e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=95e-6
mSymmetricalFirstStageStageBias12 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=418e-6
mSymmetricalFirstStageStageBias13 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=19e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias15 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
mMainBias16 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=7e-6 W=154e-6
mSymmetricalFirstStageTransconductor17 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=85e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias18 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=1e-6 W=44e-6
mSecondStage1StageBias19 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=59e-6
mSymmetricalFirstStageTransconductor20 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=85e-6
mMainBias21 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=74e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp37

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 1.09401 mW
** Area: 7383 (mu_m)^2
** Transit frequency: 3.74501 MHz
** Transit frequency with error factor: 3.74496 MHz
** Slew rate: 4.56363 V/mu_s
** Phase margin: 82.506°
** CMRR: 151 dB
** negPSRR: 51 dB
** posPSRR: 64 dB
** VoutMax: 4.51001 V
** VoutMin: 0.330001 V
** VcmMax: 3.16001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 4.86551e+07 muA
** NormalTransistorPmos: -6.69699e+06 muA
** NormalTransistorPmos: -1.40259e+07 muA
** DiodeTransistorNmos: 1.90471e+07 muA
** DiodeTransistorNmos: 1.90471e+07 muA
** NormalTransistorPmos: -3.80969e+07 muA
** NormalTransistorPmos: -3.80959e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorNmos: 4.57111e+07 muA
** NormalTransistorNmos: 4.57121e+07 muA
** NormalTransistorPmos: -4.57119e+07 muA
** NormalTransistorPmos: -4.57129e+07 muA
** NormalTransistorPmos: -4.57119e+07 muA
** NormalTransistorPmos: -4.57129e+07 muA
** NormalTransistorNmos: 4.57111e+07 muA
** NormalTransistorNmos: 4.57121e+07 muA
** DiodeTransistorNmos: 6.69601e+06 muA
** DiodeTransistorNmos: 1.40251e+07 muA
** DiodeTransistorPmos: -4.86559e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24801  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 3.91201  V
** inOutputTransconductanceComplementarySecondStage: 0.739001  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 4.15201  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.81001  V
** sourceTransconductance: 3.25701  V
** innerStageBias: 4.68401  V
** innerTransconductance: 0.150001  V
** inner: 4.71601  V
** inner: 0.150001  V


.END