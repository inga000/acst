** Name: two_stage_single_output_op_amp_58_9

.MACRO two_stage_single_output_op_amp_58_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=5e-6 W=58e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=17e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=175e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=132e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mMainBias6 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=112e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=284e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=22e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=100e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=100e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=17e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=175e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=22e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=284e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=112e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=562e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=79e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=366e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.80001e-12
.EOM two_stage_single_output_op_amp_58_9

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 2.56101 mW
** Area: 14819 (mu_m)^2
** Transit frequency: 2.54701 MHz
** Transit frequency with error factor: 2.54164 MHz
** Slew rate: 3.71774 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** VoutMax: 4.51001 V
** VoutMin: 0.700001 V
** VcmMax: 3.26001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -3.23799e+07 muA
** NormalTransistorPmos: -5.02829e+07 muA
** NormalTransistorNmos: 2.53151e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorNmos: 2.53151e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** DiodeTransistorPmos: -2.53159e+07 muA
** NormalTransistorPmos: -2.53159e+07 muA
** NormalTransistorPmos: -2.55589e+07 muA
** DiodeTransistorPmos: -2.55599e+07 muA
** NormalTransistorPmos: -1.27789e+07 muA
** NormalTransistorPmos: -1.27789e+07 muA
** NormalTransistorNmos: 3.33327e+08 muA
** DiodeTransistorNmos: 3.33326e+08 muA
** NormalTransistorPmos: -3.33326e+08 muA
** DiodeTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** DiodeTransistorNmos: 5.02821e+07 muA
** DiodeTransistorNmos: 5.02831e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.49701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.18601  V
** out: 2.5  V
** outFirstStage: 3.94801  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.24901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.97301  V
** sourceGCC1: 0.519001  V
** sourceGCC2: 0.519001  V
** sourceTransconductance: 3.29801  V
** inner: 0.555001  V
** inner: 4.24801  V


.END