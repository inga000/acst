** Name: two_stage_single_output_op_amp_66_5

.MACRO two_stage_single_output_op_amp_66_5 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=8e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
m3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=28e-6
m4 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=1e-6 W=41e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=237e-6
m6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=462e-6
m7 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=6e-6 W=40e-6
m8 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=443e-6
m9 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=62e-6
m10 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
m11 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=182e-6
m12 outVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=69e-6
m13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=62e-6
m14 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=153e-6
m15 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=153e-6
m16 out outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=462e-6
m17 outFirstStage outVoltageBiasXXpXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=268e-6
m18 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=287e-6
m19 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=287e-6
m20 FirstStageYout1 outVoltageBiasXXpXX3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=6e-6 W=268e-6
m21 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=48e-6
m22 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=48e-6
m23 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=237e-6
m24 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
m25 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_66_5

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 13.0461 mW
** Area: 9873 (mu_m)^2
** Transit frequency: 14.4661 MHz
** Transit frequency with error factor: 14.466 MHz
** Slew rate: 21.843 V/mu_s
** Phase margin: 63.5984°
** CMRR: 138 dB
** VoutMax: 3.44001 V
** VoutMin: 0.520001 V
** VcmMax: 3.32001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.17721e+07 muA
** NormalTransistorNmos: 1.80629e+08 muA
** NormalTransistorNmos: 6.76881e+07 muA
** NormalTransistorNmos: 9.98121e+07 muA
** NormalTransistorNmos: 1.50091e+08 muA
** NormalTransistorNmos: 9.98121e+07 muA
** NormalTransistorNmos: 1.50091e+08 muA
** NormalTransistorPmos: -9.98129e+07 muA
** NormalTransistorPmos: -9.98139e+07 muA
** NormalTransistorPmos: -9.98129e+07 muA
** NormalTransistorPmos: -9.98139e+07 muA
** NormalTransistorPmos: -1.00558e+08 muA
** DiodeTransistorPmos: -1.00559e+08 muA
** NormalTransistorPmos: -5.02789e+07 muA
** NormalTransistorPmos: -5.02789e+07 muA
** NormalTransistorNmos: 2.03893e+09 muA
** NormalTransistorPmos: -2.03892e+09 muA
** DiodeTransistorPmos: -2.03892e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.17729e+07 muA
** NormalTransistorPmos: -1.17739e+07 muA
** DiodeTransistorPmos: -1.80628e+08 muA
** NormalTransistorPmos: -1.80629e+08 muA
** DiodeTransistorPmos: -6.76889e+07 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.929001  V
** outInputVoltageBiasXXpXX1: 3.56401  V
** outInputVoltageBiasXXpXX2: 2.87401  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.28201  V
** outSourceVoltageBiasXXpXX2: 3.93701  V
** outVoltageBiasXXpXX3: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.60201  V
** innerTransistorStack2Load2: 4.60201  V
** out1: 4.23801  V
** sourceGCC1: 0.533001  V
** sourceGCC2: 0.533001  V
** sourceTransconductance: 3.30501  V
** inner: 4.28101  V
** inner: 3.93301  V


.END