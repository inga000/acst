.suckt  symmetrical_op_amp104 ibias in1 in2 out sourceNmos sourcePmos
mSymmetricalFirstStageLoad1 out1FirstStage out1FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mSymmetricalFirstStageLoad2 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageLoad3 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mSymmetricalFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSymmetricalFirstStageTransconductor6 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSymmetricalFirstStageTransconductor7 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1Transconductor8 out out1FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mSecondStage1Transconductor9 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias10 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos
mSecondStage1StageBias11 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias12 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor13 innerComplementarySecondStage inSourceTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mMainBias15 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp104

