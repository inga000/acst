** Name: two_stage_single_output_op_amp_34_8

.MACRO two_stage_single_output_op_amp_34_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=8e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=36e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=93e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=26e-6
m6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=13e-6
m7 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=59e-6
m8 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
m9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=55e-6
m10 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=119e-6
m11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=81e-6
m12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=81e-6
m13 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=93e-6
m14 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
m15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=36e-6
m16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=321e-6
m17 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=5e-6 W=239e-6
m18 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=197e-6
m19 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=59e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9e-12
.EOM two_stage_single_output_op_amp_34_8

** Expected Performance Values: 
** Gain: 105 dB
** Power consumption: 1.90101 mW
** Area: 10215 (mu_m)^2
** Transit frequency: 4.49801 MHz
** Transit frequency with error factor: 4.49556 MHz
** Slew rate: 4.23937 V/mu_s
** Phase margin: 60.1606°
** CMRR: 104 dB
** negPSRR: 116 dB
** posPSRR: 105 dB
** VoutMax: 4.78001 V
** VoutMin: 0.890001 V
** VcmMax: 4.39001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 1.92301e+06 muA
** NormalTransistorNmos: 2.63971e+07 muA
** NormalTransistorPmos: -1.46869e+07 muA
** DiodeTransistorPmos: -1.92859e+07 muA
** NormalTransistorPmos: -1.92859e+07 muA
** NormalTransistorPmos: -1.92859e+07 muA
** NormalTransistorNmos: 3.85691e+07 muA
** DiodeTransistorNmos: 3.85681e+07 muA
** NormalTransistorNmos: 1.92851e+07 muA
** NormalTransistorNmos: 1.92851e+07 muA
** NormalTransistorNmos: 2.88581e+08 muA
** NormalTransistorNmos: 2.8858e+08 muA
** NormalTransistorPmos: -2.8858e+08 muA
** DiodeTransistorNmos: 1.46861e+07 muA
** NormalTransistorNmos: 1.46861e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.92399e+06 muA
** DiodeTransistorPmos: -2.63979e+07 muA


** Expected Voltages: 
** ibias: 1.20201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.23201  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.21101  V
** outInputVoltageBiasXXnXX1: 1.12201  V
** outSourceVoltageBiasXXnXX1: 0.561001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.40001  V
** out1: 4.13401  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.457001  V
** inner: 0.561001  V


.END