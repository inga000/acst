** Name: two_stage_single_output_op_amp_8_9

.MACRO two_stage_single_output_op_amp_8_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=10e-6 W=37e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=304e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=87e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=24e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=8e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=10e-6 W=600e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=304e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=8e-6
mMainBias11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=59e-6
mMainBias12 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=38e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=306e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=87e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_8_9

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 3.96101 mW
** Area: 8808 (mu_m)^2
** Transit frequency: 8.25201 MHz
** Transit frequency with error factor: 8.19828 MHz
** Slew rate: 23.5058 V/mu_s
** Phase margin: 61.3065°
** CMRR: 83 dB
** negPSRR: 127 dB
** posPSRR: 81 dB
** VoutMax: 4.68001 V
** VoutMin: 0.700001 V
** VcmMax: 4.52001 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorNmos: 1.59061e+07 muA
** NormalTransistorPmos: -2.47619e+07 muA
** DiodeTransistorPmos: -8.12749e+07 muA
** NormalTransistorPmos: -8.12749e+07 muA
** NormalTransistorNmos: 1.62548e+08 muA
** NormalTransistorNmos: 8.12741e+07 muA
** NormalTransistorNmos: 8.12741e+07 muA
** NormalTransistorNmos: 5.79008e+08 muA
** DiodeTransistorNmos: 5.79008e+08 muA
** NormalTransistorPmos: -5.79007e+08 muA
** DiodeTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.59069e+07 muA


** Expected Voltages: 
** ibias: 0.583001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11001  V
** out: 2.5  V
** outFirstStage: 4.11201  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX0: 3.89401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.11201  V
** sourceTransconductance: 1.39901  V
** inner: 0.555001  V


.END