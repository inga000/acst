.suckt  complementary_op_amp12 ibias in1 in2 out sourceNmos sourcePmos
m_Complementary_MainBias_1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m_Complementary_MainBias_2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_3 FirstStageYinnerSourceLoadNmos inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m_Complementary_FirstStage_Load_4 FirstStageYinnerTransistorStack1LoadPmos outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_5 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m_Complementary_FirstStage_Load_6 FirstStageYinnerTransistorStack2LoadPmos outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_7 FirstStageYinnerSourceLoadNmos FirstStageYinnerSourceLoadNmos FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m_Complementary_FirstStage_Load_8 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_9 out FirstStageYinnerSourceLoadNmos FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m_Complementary_FirstStage_Load_10 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_11 FirstStageYsourceTransconductanceNmos ibias sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_12 FirstStageYsourceTransconductancePmos outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Transconductor_13 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_14 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_15 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m_Complementary_FirstStage_Transconductor_16 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c_Complementary_Load_Capacitor_1 out sourceNmos 
m_Complementary_MainBias_17 ibias ibias sourceNmos sourceNmos nmos
m_Complementary_MainBias_18 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_MainBias_19 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end complementary_op_amp12

