** Name: symmetrical_op_amp83

.MACRO symmetrical_op_amp83 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=8e-6
mSecondStage1StageBias2 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=150e-6
mSymmetricalFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=228e-6
mSecondStage1StageBias4 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=61e-6
mSymmetricalFirstStageLoad5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=129e-6
mSymmetricalFirstStageLoad6 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=129e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=228e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias9 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=499e-6
mSymmetricalFirstStageTransconductor10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=38e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias11 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=150e-6
mSecondStage1StageBias12 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos4 L=1e-6 W=60e-6
mSymmetricalFirstStageTransconductor13 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=38e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=171e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=171e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=456e-6
mSecondStage1Transconductor17 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=456e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp83

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 6.39601 mW
** Area: 8083 (mu_m)^2
** Transit frequency: 4.97301 MHz
** Transit frequency with error factor: 4.97263 MHz
** Slew rate: 18.4171 V/mu_s
** Phase margin: 61.3065°
** CMRR: 132 dB
** negPSRR: 46 dB
** posPSRR: 53 dB
** VoutMax: 4.25 V
** VoutMin: 0.800001 V
** VcmMax: 4.24001 V
** VcmMin: 1.74001 V


** Expected Currents: 
** NormalTransistorNmos: 6.19357e+08 muA
** DiodeTransistorPmos: -1.39709e+08 muA
** DiodeTransistorPmos: -1.39709e+08 muA
** NormalTransistorNmos: 2.79418e+08 muA
** DiodeTransistorNmos: 2.79417e+08 muA
** NormalTransistorNmos: 1.3971e+08 muA
** NormalTransistorNmos: 1.3971e+08 muA
** NormalTransistorNmos: 1.85198e+08 muA
** DiodeTransistorNmos: 1.85197e+08 muA
** NormalTransistorPmos: -1.85197e+08 muA
** NormalTransistorPmos: -1.85197e+08 muA
** NormalTransistorNmos: 1.85198e+08 muA
** NormalTransistorPmos: -1.85197e+08 muA
** NormalTransistorPmos: -1.85197e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -6.19356e+08 muA


** Expected Voltages: 
** ibias: 1.15101  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** inStageBiasComplementarySecondStage: 0.614001  V
** innerComplementarySecondStage: 1.20901  V
** out: 2.5  V
** outFirstStage: 3.83601  V
** outSourceVoltageBiasXXnXX1: 0.576001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.50301  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V
** inner: 0.574001  V


.END