** Name: two_stage_single_output_op_amp_29_10

.MACRO two_stage_single_output_op_amp_29_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
m3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=61e-6
m4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=198e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=269e-6
m6 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=501e-6
m7 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=76e-6
m8 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=302e-6
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=25e-6
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=25e-6
m11 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=241e-6
m12 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=146e-6
m13 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
m14 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=269e-6
m15 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=418e-6
m16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10.7001e-12
.EOM two_stage_single_output_op_amp_29_10

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 7.97601 mW
** Area: 8614 (mu_m)^2
** Transit frequency: 5.88801 MHz
** Transit frequency with error factor: 5.85423 MHz
** Slew rate: 12.0346 V/mu_s
** Phase margin: 60.1606°
** CMRR: 87 dB
** negPSRR: 113 dB
** posPSRR: 85 dB
** VoutMax: 4.63001 V
** VoutMin: 0.270001 V
** VcmMax: 4.66001 V
** VcmMin: 1.99001 V


** Expected Currents: 
** NormalTransistorNmos: 9.49561e+07 muA
** NormalTransistorNmos: 6.19357e+08 muA
** NormalTransistorPmos: -1.98658e+08 muA
** DiodeTransistorPmos: -1.5026e+08 muA
** NormalTransistorPmos: -1.5026e+08 muA
** NormalTransistorNmos: 3.0052e+08 muA
** NormalTransistorNmos: 3.00519e+08 muA
** NormalTransistorNmos: 1.50261e+08 muA
** NormalTransistorNmos: 1.50261e+08 muA
** NormalTransistorNmos: 3.71777e+08 muA
** NormalTransistorPmos: -3.71776e+08 muA
** NormalTransistorPmos: -3.71777e+08 muA
** DiodeTransistorNmos: 1.98659e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.49569e+07 muA
** DiodeTransistorPmos: -6.19356e+08 muA


** Expected Voltages: 
** ibias: 0.676001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.27301  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.24901  V
** outVoltageBiasXXnXX1: 0.832001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.271001  V
** out1: 4.25901  V
** sourceTransconductance: 1.34501  V
** innerTransconductance: 4.43601  V


.END