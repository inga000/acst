** Name: one_stage_single_output_op_amp61

.MACRO one_stage_single_output_op_amp61 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=7e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=173e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=16e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=52e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=121e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=121e-6
mFoldedCascodeFirstStageLoad9 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=52e-6
mMainBias10 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=186e-6
mMainBias11 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=143e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=173e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=322e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=322e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=218e-6
mFoldedCascodeFirstStageLoad17 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=25e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp61

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 2.20601 mW
** Area: 4295 (mu_m)^2
** Transit frequency: 4.85701 MHz
** Transit frequency with error factor: 4.85689 MHz
** Slew rate: 3.50001 V/mu_s
** Phase margin: 88.8085°
** CMRR: 144 dB
** VoutMax: 4.45001 V
** VoutMin: 0.740001 V
** VcmMax: 3.16001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.82761e+08 muA
** NormalTransistorNmos: 1.10081e+07 muA
** NormalTransistorNmos: 7.00621e+07 muA
** NormalTransistorNmos: 1.18701e+08 muA
** NormalTransistorNmos: 7.00591e+07 muA
** NormalTransistorNmos: 1.187e+08 muA
** DiodeTransistorPmos: -7.00609e+07 muA
** NormalTransistorPmos: -7.00599e+07 muA
** NormalTransistorPmos: -7.00609e+07 muA
** NormalTransistorPmos: -9.72789e+07 muA
** NormalTransistorPmos: -9.72799e+07 muA
** NormalTransistorPmos: -4.86389e+07 muA
** NormalTransistorPmos: -4.86389e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.8276e+08 muA
** DiodeTransistorPmos: -1.10089e+07 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.04401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40801  V
** innerTransistorStack2Load2: 4.64501  V
** out1: 4.28501  V
** sourceGCC1: 0.562001  V
** sourceGCC2: 0.562001  V
** sourceTransconductance: 3.22301  V


.END