** Name: two_stage_single_output_op_amp_29_9

.MACRO two_stage_single_output_op_amp_29_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=11e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=8e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=84e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=99e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=47e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=600e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=45e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=144e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mMainBias11 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=48e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=84e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=45e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=579e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=99e-6
mMainBias16 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=168e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.20001e-12
.EOM two_stage_single_output_op_amp_29_9

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 4.25801 mW
** Area: 8985 (mu_m)^2
** Transit frequency: 10.3681 MHz
** Transit frequency with error factor: 10.3215 MHz
** Slew rate: 21.9166 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** negPSRR: 133 dB
** posPSRR: 87 dB
** VoutMax: 4.77001 V
** VoutMin: 1.79001 V
** VcmMax: 4.61001 V
** VcmMin: 1.75 V


** Expected Currents: 
** NormalTransistorNmos: 1.53961e+07 muA
** NormalTransistorPmos: -5.39789e+07 muA
** DiodeTransistorPmos: -9.74819e+07 muA
** NormalTransistorPmos: -9.74819e+07 muA
** NormalTransistorNmos: 1.94962e+08 muA
** NormalTransistorNmos: 1.94961e+08 muA
** NormalTransistorNmos: 9.74811e+07 muA
** NormalTransistorNmos: 9.74811e+07 muA
** NormalTransistorNmos: 5.77169e+08 muA
** DiodeTransistorNmos: 5.77168e+08 muA
** NormalTransistorPmos: -5.77168e+08 muA
** DiodeTransistorNmos: 5.39781e+07 muA
** NormalTransistorNmos: 5.39781e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.53969e+07 muA


** Expected Voltages: 
** ibias: 1.21401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.10601  V
** out: 2.5  V
** outFirstStage: 4.20101  V
** outInputVoltageBiasXXnXX1: 2.20001  V
** outSourceVoltageBiasXXnXX1: 1.10001  V
** outSourceVoltageBiasXXnXX2: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.498001  V
** out1: 4.20101  V
** sourceTransconductance: 1.61301  V
** inner: 1.10001  V


.END