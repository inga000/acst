** Name: two_stage_single_output_op_amp_54_7

.MACRO two_stage_single_output_op_amp_54_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=36e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=25e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=19e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=19e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=19e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=37e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=37e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mFoldedCascodeFirstStageLoad12 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=19e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=215e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=85e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=85e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=511e-6
mFoldedCascodeFirstStageLoad17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=215e-6
mMainBias18 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=211e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=90e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.10001e-12
.EOM two_stage_single_output_op_amp_54_7

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 9.64501 mW
** Area: 8712 (mu_m)^2
** Transit frequency: 3.88701 MHz
** Transit frequency with error factor: 3.8871 MHz
** Slew rate: 3.53751 V/mu_s
** Phase margin: 60.1606°
** CMRR: 142 dB
** VoutMax: 4.25 V
** VoutMin: 0.370001 V
** VcmMax: 5.11001 V
** VcmMin: 0.940001 V


** Expected Currents: 
** NormalTransistorPmos: -8.54459e+07 muA
** NormalTransistorPmos: -3.64899e+07 muA
** NormalTransistorPmos: -2.18289e+07 muA
** NormalTransistorPmos: -3.45209e+07 muA
** NormalTransistorPmos: -2.18289e+07 muA
** NormalTransistorPmos: -3.45209e+07 muA
** NormalTransistorNmos: 2.18281e+07 muA
** NormalTransistorNmos: 2.18271e+07 muA
** NormalTransistorNmos: 2.18281e+07 muA
** NormalTransistorNmos: 2.18271e+07 muA
** NormalTransistorNmos: 2.53811e+07 muA
** NormalTransistorNmos: 1.26911e+07 muA
** NormalTransistorNmos: 1.26911e+07 muA
** NormalTransistorNmos: 1.71809e+09 muA
** NormalTransistorPmos: -1.71808e+09 muA
** DiodeTransistorNmos: 8.54451e+07 muA
** DiodeTransistorNmos: 3.64891e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.13601  V
** outVoltageBiasXXnXX1: 1.06601  V
** outVoltageBiasXXnXX2: 0.771001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.665001  V
** innerTransistorStack1Load2: 0.459001  V
** innerTransistorStack2Load2: 0.460001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.92601  V


.END