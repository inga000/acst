** Name: symmetrical_op_amp24

.MACRO symmetrical_op_amp24 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=62e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=1e-6 W=83e-6
mSecondStage1StageBias4 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSymmetricalFirstStageLoad5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=154e-6
mSymmetricalFirstStageLoad6 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=154e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=168e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=62e-6
mMainBias9 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos4 L=2e-6 W=56e-6
mSymmetricalFirstStageTransconductor10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=38e-6
mSecondStage1StageBias11 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=55e-6
mSymmetricalFirstStageTransconductor12 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=38e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=190e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=190e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=505e-6
mSecondStage1Transconductor16 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=505e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp24

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 4.32101 mW
** Area: 6401 (mu_m)^2
** Transit frequency: 5.40401 MHz
** Transit frequency with error factor: 5.40356 MHz
** Slew rate: 20.3869 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** negPSRR: 45 dB
** posPSRR: 53 dB
** VoutMax: 4.25 V
** VoutMin: 0.810001 V
** VcmMax: 4.24001 V
** VcmMin: 1.23001 V


** Expected Currents: 
** NormalTransistorNmos: 1.1053e+08 muA
** DiodeTransistorPmos: -1.66785e+08 muA
** DiodeTransistorPmos: -1.66785e+08 muA
** NormalTransistorNmos: 3.3357e+08 muA
** NormalTransistorNmos: 1.66786e+08 muA
** NormalTransistorNmos: 1.66786e+08 muA
** NormalTransistorNmos: 2.05098e+08 muA
** NormalTransistorNmos: 2.05097e+08 muA
** NormalTransistorPmos: -2.05097e+08 muA
** NormalTransistorPmos: -2.05098e+08 muA
** DiodeTransistorNmos: 2.05098e+08 muA
** DiodeTransistorNmos: 2.05097e+08 muA
** NormalTransistorPmos: -2.05097e+08 muA
** NormalTransistorPmos: -2.05098e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.10529e+08 muA


** Expected Voltages: 
** ibias: 0.622001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceStageBiasComplementarySecondStage: 0.602001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 1.17701  V
** out: 2.5  V
** outFirstStage: 3.83601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.49001  V
** innerStageBias: 0.562001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END