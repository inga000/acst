** Name: two_stage_single_output_op_amp_5_5

.MACRO two_stage_single_output_op_amp_5_5 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=40e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=17e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=26e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=229e-6
m6 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=134e-6
m7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=122e-6
m8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=122e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=598e-6
m10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=134e-6
m11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=102e-6
m12 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=279e-6
m13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=597e-6
m14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
m15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=369e-6
m16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=229e-6
m17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=279e-6
m18 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_5_5

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 12.2361 mW
** Area: 4971 (mu_m)^2
** Transit frequency: 28.6431 MHz
** Transit frequency with error factor: 28.5987 MHz
** Slew rate: 46.2791 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 100 dB
** posPSRR: 125 dB
** VoutMax: 3.28001 V
** VoutMin: 0.160001 V
** VcmMax: 3.88001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorNmos: 1.56789e+08 muA
** NormalTransistorPmos: -2.58139e+07 muA
** NormalTransistorPmos: -3.39016e+08 muA
** NormalTransistorNmos: 2.75201e+08 muA
** NormalTransistorNmos: 2.752e+08 muA
** NormalTransistorNmos: 2.75201e+08 muA
** NormalTransistorNmos: 2.752e+08 muA
** NormalTransistorPmos: -5.50401e+08 muA
** NormalTransistorPmos: -2.752e+08 muA
** NormalTransistorPmos: -2.752e+08 muA
** NormalTransistorNmos: 1.35526e+09 muA
** NormalTransistorPmos: -1.35525e+09 muA
** DiodeTransistorPmos: -1.35525e+09 muA
** DiodeTransistorNmos: 2.58131e+07 muA
** DiodeTransistorNmos: 3.39017e+08 muA
** DiodeTransistorPmos: -1.56788e+08 muA
** NormalTransistorPmos: -1.56788e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.723001  V
** out: 2.5  V
** outFirstStage: 0.568001  V
** outInputVoltageBiasXXpXX1: 2.71601  V
** outSourceVoltageBiasXXpXX1: 3.85801  V
** outVoltageBiasXXnXX0: 0.829001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.568001  V
** innerTransistorStack1Load1: 0.163001  V
** innerTransistorStack2Load1: 0.163001  V
** sourceTransconductance: 3.39501  V
** inner: 3.85801  V


.END