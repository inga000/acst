** Name: two_stage_single_output_op_amp_24_2

.MACRO two_stage_single_output_op_amp_24_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=19e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=56e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=19e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=140e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=330e-6
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=23e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=69e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=69e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=168e-6
mSecondStage1Transconductor10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=168e-6
mSimpleFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=23e-6
mMainBias12 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=71e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=291e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=330e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=140e-6
mMainBias16 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=269e-6
mSecondStage1StageBias17 out ibias sourcePmos sourcePmos pmos4 L=4e-6 W=600e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=291e-6
mMainBias19 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=55e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.60001e-12
.EOM two_stage_single_output_op_amp_24_2

** Expected Performance Values: 
** Gain: 104 dB
** Power consumption: 3.19201 mW
** Area: 12705 (mu_m)^2
** Transit frequency: 7.03101 MHz
** Transit frequency with error factor: 7.02465 MHz
** Slew rate: 9.06725 V/mu_s
** Phase margin: 60.1606°
** CMRR: 104 dB
** negPSRR: 105 dB
** posPSRR: 168 dB
** VoutMax: 4.66001 V
** VoutMin: 0.300001 V
** VcmMax: 3.12001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.76671e+07 muA
** NormalTransistorPmos: -2.93699e+07 muA
** NormalTransistorPmos: -1.43319e+08 muA
** NormalTransistorNmos: 4.38101e+07 muA
** NormalTransistorNmos: 4.38091e+07 muA
** NormalTransistorNmos: 4.38101e+07 muA
** NormalTransistorNmos: 4.38091e+07 muA
** NormalTransistorPmos: -8.76229e+07 muA
** DiodeTransistorPmos: -8.76239e+07 muA
** NormalTransistorPmos: -4.38109e+07 muA
** NormalTransistorPmos: -4.38109e+07 muA
** NormalTransistorNmos: 3.20403e+08 muA
** NormalTransistorNmos: 3.20402e+08 muA
** NormalTransistorPmos: -3.20402e+08 muA
** DiodeTransistorNmos: 2.93691e+07 muA
** DiodeTransistorNmos: 1.4332e+08 muA
** DiodeTransistorPmos: -3.76679e+07 muA
** NormalTransistorPmos: -3.76679e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.09201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.32601  V
** outSourceVoltageBiasXXpXX1: 4.16301  V
** outVoltageBiasXXnXX0: 0.563001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.26901  V
** innerTransconductance: 0.150001  V
** inner: 4.16301  V


.END