** Name: two_stage_single_output_op_amp_58_12

.MACRO two_stage_single_output_op_amp_58_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=6e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=491e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
mMainBias6 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=236e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=195e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=43e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=43e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=6e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=491e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=195e-6
mMainBias15 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=482e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=482e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=236e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=547e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias21 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=33e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=585e-6
mFoldedCascodeFirstStageLoad23 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
mMainBias24 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14e-12
.EOM two_stage_single_output_op_amp_58_12

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 10.9021 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 8.12701 MHz
** Transit frequency with error factor: 8.11448 MHz
** Slew rate: 11.9981 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** VoutMax: 4.25 V
** VoutMin: 1.14001 V
** VcmMax: 3.06001 V
** VcmMin: -0.0799999 V


** Expected Currents: 
** NormalTransistorNmos: 1.00565e+08 muA
** NormalTransistorPmos: -1.72349e+07 muA
** NormalTransistorPmos: -3.28599e+07 muA
** NormalTransistorNmos: 1.68649e+08 muA
** NormalTransistorNmos: 2.88286e+08 muA
** NormalTransistorNmos: 1.68649e+08 muA
** NormalTransistorNmos: 2.88286e+08 muA
** DiodeTransistorPmos: -1.68648e+08 muA
** NormalTransistorPmos: -1.68648e+08 muA
** NormalTransistorPmos: -2.39275e+08 muA
** DiodeTransistorPmos: -2.39274e+08 muA
** NormalTransistorPmos: -1.19637e+08 muA
** NormalTransistorPmos: -1.19637e+08 muA
** NormalTransistorNmos: 1.43327e+09 muA
** DiodeTransistorNmos: 1.43327e+09 muA
** NormalTransistorPmos: -1.43326e+09 muA
** NormalTransistorPmos: -1.43326e+09 muA
** DiodeTransistorNmos: 1.72341e+07 muA
** NormalTransistorNmos: 1.72331e+07 muA
** DiodeTransistorNmos: 3.28591e+07 muA
** DiodeTransistorNmos: 3.28581e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.00564e+08 muA


** Expected Voltages: 
** ibias: 3.39601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.77601  V
** out: 2.5  V
** outFirstStage: 4.05501  V
** outInputVoltageBiasXXnXX1: 1.55001  V
** outSourceVoltageBiasXXnXX1: 0.775001  V
** outSourceVoltageBiasXXnXX2: 0.890001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.04401  V
** sourceGCC1: 1.19601  V
** sourceGCC2: 1.19601  V
** sourceTransconductance: 3.39601  V
** innerTransconductance: 4.61901  V
** inner: 0.775001  V
** inner: 4.19601  V


.END