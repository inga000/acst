** Name: symmetrical_op_amp24

.MACRO symmetrical_op_amp24 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
m2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=92e-6
m3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=1e-6 W=179e-6
m4 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
m6 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
m7 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos4 L=2e-6 W=61e-6
m8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=43e-6
m9 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=156e-6
m10 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=43e-6
m11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=461e-6
m12 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=92e-6
m13 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=599e-6
m14 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
m15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=59e-6
m16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=59e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp24

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 7.82201 mW
** Area: 3117 (mu_m)^2
** Transit frequency: 16.9371 MHz
** Transit frequency with error factor: 16.9373 MHz
** Slew rate: 33.9778 V/mu_s
** Phase margin: 82.506°
** CMRR: 137 dB
** negPSRR: 51 dB
** posPSRR: 57 dB
** VoutMax: 4.25 V
** VoutMin: 0.770001 V
** VcmMax: 4.27001 V
** VcmMin: 0.930001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** DiodeTransistorPmos: -3.83878e+08 muA
** DiodeTransistorPmos: -3.83878e+08 muA
** NormalTransistorNmos: 7.67756e+08 muA
** NormalTransistorNmos: 3.83879e+08 muA
** NormalTransistorNmos: 3.83879e+08 muA
** NormalTransistorNmos: 3.42575e+08 muA
** NormalTransistorNmos: 3.42574e+08 muA
** NormalTransistorPmos: -3.42574e+08 muA
** NormalTransistorPmos: -3.42575e+08 muA
** DiodeTransistorNmos: 3.42575e+08 muA
** DiodeTransistorNmos: 3.42574e+08 muA
** NormalTransistorPmos: -3.42574e+08 muA
** NormalTransistorPmos: -3.42575e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceStageBiasComplementarySecondStage: 0.614001  V
** inSourceTransconductanceComplementarySecondStage: 3.86401  V
** innerComplementarySecondStage: 1.16901  V
** out: 2.5  V
** outFirstStage: 3.86401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.76901  V
** innerStageBias: 0.603001  V
** innerTransconductance: 4.42801  V
** inner: 4.42801  V


.END