.suckt  two_stage_fully_differential_op_amp_32_7 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m5 outFeedback outFeedback sourceNmos sourceNmos nmos
m6 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m7 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m8 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m9 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m14 out1FirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m15 FirstStageYinnerTransistorStack1Load1 outFeedback sourceNmos sourceNmos nmos
m16 out2FirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m17 FirstStageYinnerTransistorStack2Load1 outFeedback sourceNmos sourceNmos nmos
m18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m19 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m20 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m21 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m22 out1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m23 out1 out1FirstStage sourcePmos sourcePmos pmos
m24 out2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m25 out2 out2FirstStage sourcePmos sourcePmos pmos
m26 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m27 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m28 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m29 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m30 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m31 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_32_7

