** Name: two_stage_single_output_op_amp_44_2

.MACRO two_stage_single_output_op_amp_44_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=6e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=271e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=30e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=49e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=137e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=137e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=282e-6
mSecondStage1Transconductor9 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=205e-6
mFoldedCascodeFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=49e-6
mFoldedCascodeFirstStageLoad11 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=9e-6 W=271e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=25e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=25e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=162e-6
mMainBias15 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=13e-6
mSecondStage1StageBias16 out ibias sourcePmos sourcePmos pmos4 L=4e-6 W=597e-6
mFoldedCascodeFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=9e-6 W=286e-6
mMainBias18 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=96e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_44_2

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 1.95201 mW
** Area: 14967 (mu_m)^2
** Transit frequency: 2.72701 MHz
** Transit frequency with error factor: 2.72657 MHz
** Slew rate: 8.20095 V/mu_s
** Phase margin: 69.328°
** CMRR: 126 dB
** VoutMax: 4.73001 V
** VoutMin: 0.400001 V
** VcmMax: 3.46001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -3.21069e+07 muA
** NormalTransistorPmos: -4.31799e+06 muA
** NormalTransistorNmos: 3.84181e+07 muA
** NormalTransistorNmos: 6.58611e+07 muA
** NormalTransistorNmos: 3.84151e+07 muA
** NormalTransistorNmos: 6.58561e+07 muA
** NormalTransistorPmos: -3.84169e+07 muA
** NormalTransistorPmos: -3.84159e+07 muA
** DiodeTransistorPmos: -3.84169e+07 muA
** NormalTransistorPmos: -5.48829e+07 muA
** NormalTransistorPmos: -2.74419e+07 muA
** NormalTransistorPmos: -2.74419e+07 muA
** NormalTransistorNmos: 2.02257e+08 muA
** NormalTransistorNmos: 2.02256e+08 muA
** NormalTransistorPmos: -2.02256e+08 muA
** DiodeTransistorNmos: 3.21061e+07 muA
** DiodeTransistorNmos: 4.31701e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.16201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.565001  V
** outVoltageBiasXXnXX1: 0.970001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.16801  V
** out1: 3.34301  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.76201  V
** innerTransconductance: 0.323001  V


.END