** Name: two_stage_single_output_op_amp_24_1

.MACRO two_stage_single_output_op_amp_24_1 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=170e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=59e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=33e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=278e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=75e-6
m6 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=410e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=80e-6
m8 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=244e-6
m9 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=8e-6 W=80e-6
m10 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m11 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m12 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=527e-6
m13 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=367e-6
m14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=130e-6
m15 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=111e-6
m16 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=130e-6
m17 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=75e-6
m18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=278e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_24_1

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 2.53801 mW
** Area: 13119 (mu_m)^2
** Transit frequency: 2.58601 MHz
** Transit frequency with error factor: 2.58245 MHz
** Slew rate: 3.8126 V/mu_s
** Phase margin: 60.1606°
** CMRR: 102 dB
** negPSRR: 103 dB
** posPSRR: 197 dB
** VoutMax: 4.82001 V
** VoutMin: 0.150001 V
** VcmMax: 3.28001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.43319e+08 muA
** NormalTransistorPmos: -3.42859e+07 muA
** NormalTransistorPmos: -1.60291e+08 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorPmos: -3.80929e+07 muA
** DiodeTransistorPmos: -3.80939e+07 muA
** NormalTransistorPmos: -1.90469e+07 muA
** NormalTransistorPmos: -1.90469e+07 muA
** NormalTransistorNmos: 1.11558e+08 muA
** NormalTransistorPmos: -1.11557e+08 muA
** DiodeTransistorNmos: 3.42851e+07 muA
** DiodeTransistorNmos: 1.60292e+08 muA
** DiodeTransistorPmos: -1.43318e+08 muA
** NormalTransistorPmos: -1.43319e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.53401  V
** outSourceVoltageBiasXXpXX1: 4.26701  V
** outVoltageBiasXXnXX0: 0.654001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.31901  V
** inner: 4.26701  V


.END