** Name: one_stage_single_output_op_amp65

.MACRO one_stage_single_output_op_amp65 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=10e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=126e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=376e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=376e-6
mFoldedCascodeFirstStageLoad8 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=126e-6
mMainBias9 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=62e-6
mMainBias10 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=26e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=115e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=108e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=108e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=413e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=317e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=317e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=443e-6
mFoldedCascodeFirstStageLoad18 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=413e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp65

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 2.79901 mW
** Area: 7516 (mu_m)^2
** Transit frequency: 7.68001 MHz
** Transit frequency with error factor: 7.68033 MHz
** Slew rate: 8.0885 V/mu_s
** Phase margin: 86.5167°
** CMRR: 139 dB
** VoutMax: 4.5 V
** VoutMin: 0.770001 V
** VcmMax: 3.21001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.06121e+07 muA
** NormalTransistorNmos: 1.73471e+07 muA
** NormalTransistorNmos: 1.62718e+08 muA
** NormalTransistorNmos: 2.459e+08 muA
** NormalTransistorNmos: 1.62718e+08 muA
** NormalTransistorNmos: 2.459e+08 muA
** NormalTransistorPmos: -1.62717e+08 muA
** NormalTransistorPmos: -1.62718e+08 muA
** NormalTransistorPmos: -1.62717e+08 muA
** NormalTransistorPmos: -1.62718e+08 muA
** NormalTransistorPmos: -1.66366e+08 muA
** NormalTransistorPmos: -1.66367e+08 muA
** NormalTransistorPmos: -8.31829e+07 muA
** NormalTransistorPmos: -8.31829e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -4.06129e+07 muA
** DiodeTransistorPmos: -1.73479e+07 muA


** Expected Voltages: 
** ibias: 1.15101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.15101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.45401  V
** innerTransistorStack1Load2: 4.45901  V
** innerTransistorStack2Load2: 4.45901  V
** out1: 4.14501  V
** sourceGCC1: 0.531001  V
** sourceGCC2: 0.531001  V
** sourceTransconductance: 3.23501  V


.END