** Name: one_stage_single_output_op_amp44

.MACRO one_stage_single_output_op_amp44 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=33e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=19e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=10e-6 W=83e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=144e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=129e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=129e-6
mFoldedCascodeFirstStageLoad8 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=144e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=64e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=64e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=10e-6 W=594e-6
mMainBias13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=10e-6 W=130e-6
mFoldedCascodeFirstStageLoad14 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp44

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 1.24201 mW
** Area: 10640 (mu_m)^2
** Transit frequency: 3.23401 MHz
** Transit frequency with error factor: 3.23411 MHz
** Slew rate: 3.5 V/mu_s
** Phase margin: 86.5167°
** CMRR: 130 dB
** VoutMax: 3.36001 V
** VoutMin: 0.75 V
** VcmMax: 4 V
** VcmMin: -0.369999 V


** Expected Currents: 
** NormalTransistorPmos: -1.57149e+07 muA
** NormalTransistorNmos: 7.01311e+07 muA
** NormalTransistorNmos: 1.06371e+08 muA
** NormalTransistorNmos: 7.01281e+07 muA
** NormalTransistorNmos: 1.06368e+08 muA
** NormalTransistorPmos: -7.01299e+07 muA
** NormalTransistorPmos: -7.01289e+07 muA
** DiodeTransistorPmos: -7.01299e+07 muA
** NormalTransistorPmos: -7.24799e+07 muA
** NormalTransistorPmos: -3.62399e+07 muA
** NormalTransistorPmos: -3.62399e+07 muA
** DiodeTransistorNmos: 1.57141e+07 muA
** DiodeTransistorNmos: 1.57131e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.15701  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.602001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 3.99101  V
** out1: 2.79801  V
** sourceGCC1: 0.600001  V
** sourceGCC2: 0.600001  V
** sourceTransconductance: 3.24201  V


.END