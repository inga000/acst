** Name: two_stage_single_output_op_amp_44_9

.MACRO two_stage_single_output_op_amp_44_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=41e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=39e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=562e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=385e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=38e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=32e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=107e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=107e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=562e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=32e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=385e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=160e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=160e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=598e-6
mMainBias17 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=577e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=414e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=3e-6 W=162e-6
mMainBias20 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=547e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.7001e-12
.EOM two_stage_single_output_op_amp_44_9

** Expected Performance Values: 
** Gain: 115 dB
** Power consumption: 14.4501 mW
** Area: 13655 (mu_m)^2
** Transit frequency: 8.15701 MHz
** Transit frequency with error factor: 8.15704 MHz
** Slew rate: 14.5039 V/mu_s
** Phase margin: 60.1606°
** CMRR: 126 dB
** VoutMax: 4.25 V
** VoutMin: 1 V
** VcmMax: 3.91001 V
** VcmMin: -0.289999 V


** Expected Currents: 
** NormalTransistorPmos: -1.45755e+08 muA
** NormalTransistorPmos: -1.51139e+08 muA
** NormalTransistorNmos: 1.55957e+08 muA
** NormalTransistorNmos: 2.35629e+08 muA
** NormalTransistorNmos: 1.55956e+08 muA
** NormalTransistorNmos: 2.35628e+08 muA
** NormalTransistorPmos: -1.55956e+08 muA
** NormalTransistorPmos: -1.55955e+08 muA
** DiodeTransistorPmos: -1.55956e+08 muA
** NormalTransistorPmos: -1.59345e+08 muA
** NormalTransistorPmos: -7.96729e+07 muA
** NormalTransistorPmos: -7.96729e+07 muA
** NormalTransistorNmos: 2.10176e+09 muA
** DiodeTransistorNmos: 2.10176e+09 muA
** NormalTransistorPmos: -2.10175e+09 muA
** DiodeTransistorNmos: 1.45756e+08 muA
** NormalTransistorNmos: 1.45755e+08 muA
** DiodeTransistorNmos: 1.5114e+08 muA
** DiodeTransistorNmos: 1.51139e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.44801  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.40201  V
** outSourceVoltageBiasXXnXX1: 0.701001  V
** outSourceVoltageBiasXXnXX2: 0.683001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.28601  V
** out1: 3.32201  V
** sourceGCC1: 0.626001  V
** sourceGCC2: 0.626001  V
** sourceTransconductance: 3.35201  V
** inner: 0.699001  V


.END