** Name: two_stage_single_output_op_amp_8_10

.MACRO two_stage_single_output_op_amp_8_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=169e-6
mSecondStage1StageBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSimpleFirstStageTransconductor4 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=104e-6
mSimpleFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=86e-6
mSecondStage1StageBias6 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mSimpleFirstStageTransconductor7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=104e-6
mMainBias8 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=135e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=548e-6
mSecondStage1Transconductor10 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=589e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=169e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.4001e-12
.EOM two_stage_single_output_op_amp_8_10

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 3.42601 mW
** Area: 7080 (mu_m)^2
** Transit frequency: 6.31801 MHz
** Transit frequency with error factor: 6.31072 MHz
** Slew rate: 6.15939 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 166 dB
** posPSRR: 98 dB
** VoutMax: 4.56001 V
** VoutMin: 0.200001 V
** VcmMax: 4.62001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorNmos: 1.11687e+08 muA
** DiodeTransistorPmos: -3.53229e+07 muA
** NormalTransistorPmos: -3.53229e+07 muA
** NormalTransistorNmos: 7.06441e+07 muA
** NormalTransistorNmos: 3.53221e+07 muA
** NormalTransistorNmos: 3.53221e+07 muA
** NormalTransistorNmos: 4.92866e+08 muA
** NormalTransistorPmos: -4.92865e+08 muA
** NormalTransistorPmos: -4.92866e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.11686e+08 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.21101  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.21901  V
** sourceTransconductance: 1.94001  V
** innerTransconductance: 4.46601  V


.END