** Name: one_stage_single_output_op_amp82

.MACRO one_stage_single_output_op_amp82 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=8e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=149e-6
m3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=20e-6
m5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=42e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m7 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=49e-6
m8 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=20e-6
m9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=66e-6
m11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=66e-6
m12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=149e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
m14 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=373e-6
m15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=373e-6
m16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=45e-6
m17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=45e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp82

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 2.78501 mW
** Area: 2522 (mu_m)^2
** Transit frequency: 8.02101 MHz
** Transit frequency with error factor: 8.02068 MHz
** Slew rate: 7.53843 V/mu_s
** Phase margin: 87.0896°
** CMRR: 140 dB
** VoutMax: 3.73001 V
** VoutMin: 1.43001 V
** VcmMax: 4.85001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorNmos: 6.05001e+07 muA
** NormalTransistorPmos: -1.51487e+08 muA
** NormalTransistorPmos: -2.43274e+08 muA
** NormalTransistorPmos: -1.51487e+08 muA
** NormalTransistorPmos: -2.43274e+08 muA
** DiodeTransistorNmos: 1.51488e+08 muA
** NormalTransistorNmos: 1.51487e+08 muA
** NormalTransistorNmos: 1.51488e+08 muA
** DiodeTransistorNmos: 1.51487e+08 muA
** NormalTransistorNmos: 1.83574e+08 muA
** DiodeTransistorNmos: 1.83575e+08 muA
** NormalTransistorNmos: 9.17861e+07 muA
** NormalTransistorNmos: 9.17861e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -6.05009e+07 muA
** DiodeTransistorPmos: -6.05e+07 muA


** Expected Voltages: 
** ibias: 1.22801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.615001  V
** outSourceVoltageBiasXXpXX1: 3.88401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 1.13301  V
** innerTransistorStack2Load2: 1.13501  V
** out1: 1.83801  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.91301  V
** inner: 0.612001  V


.END