.suckt  two_stage_fully_differential_op_amp_37_2 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m5 outFeedback outFeedback sourceNmos sourceNmos nmos
m6 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m7 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m8 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m9 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m10 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m12 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m13 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m14 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m15 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m16 out1FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m17 FirstStageYinnerTransistorStack1Load2 ibias sourcePmos sourcePmos pmos
m18 out2FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m19 FirstStageYinnerTransistorStack2Load2 ibias sourcePmos sourcePmos pmos
m20 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m21 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
m22 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m23 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m24 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m25 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m26 out1 ibias sourcePmos sourcePmos pmos
m27 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m28 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m29 out2 ibias sourcePmos sourcePmos pmos
m30 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m31 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m32 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m33 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_37_2

