** Name: two_stage_single_output_op_amp_78_2

.MACRO two_stage_single_output_op_amp_78_2 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=5e-6 W=44e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=25e-6
mMainBias3 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=15e-6
mSecondStage1StageBias4 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=36e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=78e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=213e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=5e-6 W=44e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=11e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=11e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=36e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=34e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSecondStage1Transconductor14 out inputVoltageBiasXXnXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=452e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=25e-6
mMainBias16 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=594e-6
mMainBias17 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=375e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=37e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mFoldedCascodeFirstStageLoad20 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mMainBias21 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=306e-6
mSecondStage1StageBias22 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=374e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=37e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_78_2

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 7.46601 mW
** Area: 6266 (mu_m)^2
** Transit frequency: 3.30001 MHz
** Transit frequency with error factor: 3.29988 MHz
** Slew rate: 3.71127 V/mu_s
** Phase margin: 63.0254°
** CMRR: 137 dB
** VoutMax: 4.75 V
** VoutMin: 0.700001 V
** VcmMax: 5.15001 V
** VcmMin: 1.37001 V


** Expected Currents: 
** NormalTransistorNmos: 3.95982e+08 muA
** NormalTransistorNmos: 2.46099e+08 muA
** NormalTransistorPmos: -3.53549e+08 muA
** NormalTransistorPmos: -1.67609e+07 muA
** NormalTransistorPmos: -2.85329e+07 muA
** NormalTransistorPmos: -1.67609e+07 muA
** NormalTransistorPmos: -2.85329e+07 muA
** DiodeTransistorNmos: 1.67601e+07 muA
** DiodeTransistorNmos: 1.67611e+07 muA
** NormalTransistorNmos: 1.67601e+07 muA
** NormalTransistorNmos: 1.67611e+07 muA
** NormalTransistorNmos: 2.35431e+07 muA
** DiodeTransistorNmos: 2.35441e+07 muA
** NormalTransistorNmos: 1.17711e+07 muA
** NormalTransistorNmos: 1.17711e+07 muA
** NormalTransistorNmos: 4.30447e+08 muA
** NormalTransistorNmos: 4.30446e+08 muA
** NormalTransistorPmos: -4.30446e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 3.5355e+08 muA
** DiodeTransistorPmos: -3.95981e+08 muA
** DiodeTransistorPmos: -2.46098e+08 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.10301  V
** out: 2.5  V
** outFirstStage: 0.953001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.18301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.554001  V
** out1: 1.15801  V
** sourceGCC1: 4.47501  V
** sourceGCC2: 4.47501  V
** sourceTransconductance: 1.84301  V
** innerTransconductance: 0.548001  V
** inner: 0.556001  V


.END