** Name: two_stage_single_output_op_amp_40_8

.MACRO two_stage_single_output_op_amp_40_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=7e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=536e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=54e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=54e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=54e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=486e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=49e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=54e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=536e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mSecondStage1StageBias13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=211e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=49e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=54e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=451e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=54e-6
mMainBias18 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=382e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_40_8

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 8.51101 mW
** Area: 14714 (mu_m)^2
** Transit frequency: 5.36501 MHz
** Transit frequency with error factor: 5.36166 MHz
** Slew rate: 5.05607 V/mu_s
** Phase margin: 60.1606°
** CMRR: 106 dB
** negPSRR: 109 dB
** posPSRR: 100 dB
** VoutMax: 4.61001 V
** VoutMin: 0.820001 V
** VcmMax: 3.90001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorNmos: 5.90216e+08 muA
** NormalTransistorPmos: -4.54848e+08 muA
** DiodeTransistorPmos: -2.33329e+07 muA
** NormalTransistorPmos: -2.33339e+07 muA
** NormalTransistorPmos: -2.33329e+07 muA
** DiodeTransistorPmos: -2.33339e+07 muA
** NormalTransistorNmos: 4.66631e+07 muA
** DiodeTransistorNmos: 4.66621e+07 muA
** NormalTransistorNmos: 2.33321e+07 muA
** NormalTransistorNmos: 2.33321e+07 muA
** NormalTransistorNmos: 6.00478e+08 muA
** NormalTransistorNmos: 6.00477e+08 muA
** NormalTransistorPmos: -6.00477e+08 muA
** DiodeTransistorNmos: 4.54849e+08 muA
** NormalTransistorNmos: 4.54849e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.90215e+08 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.85601  V
** out: 2.5  V
** outFirstStage: 4.04901  V
** outInputVoltageBiasXXnXX1: 1.26001  V
** outSourceVoltageBiasXXnXX1: 0.630001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.28001  V
** innerTransistorStack1Load1: 4.27801  V
** out1: 3.49501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.481001  V
** inner: 0.630001  V


.END