** Name: two_stage_single_output_op_amp_50_10

.MACRO two_stage_single_output_op_amp_50_10 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=199e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=9e-6
mMainBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=97e-6
mFoldedCascodeFirstStageTransconductor5 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=21e-6
mFoldedCascodeFirstStageTransconductor6 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=21e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=177e-6
mSecondStage1StageBias8 out ibias sourceNmos sourceNmos nmos4 L=7e-6 W=589e-6
mFoldedCascodeFirstStageLoad9 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=199e-6
mMainBias10 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=92e-6
mMainBias11 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=40e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=222e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=548e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=548e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=530e-6
mSecondStage1Transconductor16 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=600e-6
mFoldedCascodeFirstStageLoad17 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=222e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.2001e-12
.EOM two_stage_single_output_op_amp_50_10

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 6.50401 mW
** Area: 14818 (mu_m)^2
** Transit frequency: 3.69701 MHz
** Transit frequency with error factor: 3.68921 MHz
** Slew rate: 13.5523 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** VoutMax: 4.25 V
** VoutMin: 0.300001 V
** VcmMax: 5.25 V
** VcmMin: 1.45001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorNmos: 4.42631e+07 muA
** NormalTransistorPmos: -1.53155e+08 muA
** NormalTransistorPmos: -2.5007e+08 muA
** NormalTransistorPmos: -1.53155e+08 muA
** NormalTransistorPmos: -2.5007e+08 muA
** DiodeTransistorNmos: 1.53156e+08 muA
** NormalTransistorNmos: 1.53156e+08 muA
** NormalTransistorNmos: 1.93828e+08 muA
** NormalTransistorNmos: 9.69141e+07 muA
** NormalTransistorNmos: 9.69141e+07 muA
** NormalTransistorNmos: 6.44792e+08 muA
** NormalTransistorPmos: -6.44791e+08 muA
** NormalTransistorPmos: -6.44792e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -4.42639e+07 muA


** Expected Voltages: 
** ibias: 0.707001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.17401  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.27701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.618001  V
** sourceGCC1: 4.64101  V
** sourceGCC2: 4.64101  V
** sourceTransconductance: 1.35301  V
** innerTransconductance: 4.73801  V


.END