.suckt  complementary_op_amp1 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 FirstStageYinnerOutputLoadPmos FirstStageYinnerOutputLoadPmos FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos pmos
m3 FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m4 out FirstStageYinnerOutputLoadPmos FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m5 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m6 FirstStageYinnerOutputLoadPmos FirstStageYinnerOutputLoadPmos FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m7 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos sourceNmos sourceNmos nmos
m8 out FirstStageYinnerOutputLoadPmos FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m9 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack1LoadNmos sourceNmos sourceNmos nmos
m10 FirstStageYsourceTransconductanceNmos outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m11 FirstStageYsourceTransconductancePmos ibias sourcePmos sourcePmos pmos
m12 FirstStageYinnerSourceLoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m13 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m14 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m15 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c1 out sourceNmos 
m16 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m17 ibias ibias sourcePmos sourcePmos pmos
.end complementary_op_amp1

