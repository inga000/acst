.suckt  symmetrical_op_amp119 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_MainBias_1 out2FirstStage ibias sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Load_2 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m_Symmetrical_FirstStage_Load_3 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_4 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_Symmetrical_FirstStage_Load_5 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_StageBias_6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Transconductor_7 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_Symmetrical_FirstStage_Transconductor_8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_StageBias_9 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos
m_Symmetrical_SecondStage1_StageBias_10 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_Transconductor_11 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m_Symmetrical_SecondStage1_Transconductor_12 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_13 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_14 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_15 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_MainBias_17 ibias ibias sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_18 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos
.end symmetrical_op_amp119

