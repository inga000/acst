** Name: two_stage_single_output_op_amp_9_8

.MACRO two_stage_single_output_op_amp_9_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=39e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=20e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=9e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=14e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=237e-6
mSecondStage1StageBias8 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=225e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=9e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mSimpleFirstStageLoad11 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=39e-6
mMainBias12 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=51e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=138e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=9e-6 W=114e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5e-12
.EOM two_stage_single_output_op_amp_9_8

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 2.80301 mW
** Area: 5270 (mu_m)^2
** Transit frequency: 2.88901 MHz
** Transit frequency with error factor: 2.88539 MHz
** Slew rate: 5.44838 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 97 dB
** posPSRR: 88 dB
** VoutMax: 4.25 V
** VoutMin: 0.690001 V
** VcmMax: 4.17001 V
** VcmMin: 1.05001 V


** Expected Currents: 
** NormalTransistorNmos: 1.59741e+07 muA
** NormalTransistorPmos: -4.00199e+07 muA
** NormalTransistorPmos: -1.37249e+07 muA
** NormalTransistorPmos: -1.37249e+07 muA
** DiodeTransistorPmos: -1.37249e+07 muA
** NormalTransistorNmos: 2.74491e+07 muA
** NormalTransistorNmos: 1.37241e+07 muA
** NormalTransistorNmos: 1.37241e+07 muA
** NormalTransistorNmos: 4.67056e+08 muA
** NormalTransistorNmos: 4.67055e+08 muA
** NormalTransistorPmos: -4.67055e+08 muA
** DiodeTransistorNmos: 4.00191e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.59749e+07 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.09601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 3.84101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.01501  V
** out1: 3.20501  V
** sourceTransconductance: 1.79401  V
** innerStageBias: 0.342001  V


.END