.suckt  two_stage_fully_differential_op_amp_49_8 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m3 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m4 outFeedback outFeedback sourcePmos sourcePmos pmos
m5 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m6 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m7 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m8 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m9 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m10 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m11 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m12 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m13 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m14 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m15 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m16 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m17 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias nmos
m18 SecondStage1YinnerStageBias ibias sourceNmos sourceNmos nmos
m19 out1 out1FirstStage sourcePmos sourcePmos pmos
m20 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias nmos
m21 SecondStage2YinnerStageBias ibias sourceNmos sourceNmos nmos
m22 out2 out2FirstStage sourcePmos sourcePmos pmos
m23 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m24 ibias ibias sourceNmos sourceNmos nmos
m25 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_49_8

