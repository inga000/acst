** Name: symmetrical_op_amp94

.MACRO symmetrical_op_amp94 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m2 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=34e-6
m3 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
m4 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=11e-6
m5 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=19e-6
m6 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=1e-6 W=47e-6
m7 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=47e-6
m8 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=19e-6
m9 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
m10 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
m11 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=172e-6
m12 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=172e-6
m13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=124e-6
m14 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=203e-6
m15 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=124e-6
m16 out2FirstStage ibias sourcePmos sourcePmos pmos4 L=4e-6 W=281e-6
m17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=299e-6
m18 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp94

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 2.06101 mW
** Area: 5858 (mu_m)^2
** Transit frequency: 5.00101 MHz
** Transit frequency with error factor: 5.00113 MHz
** Slew rate: 10.9886 V/mu_s
** Phase margin: 79.0682°
** CMRR: 147 dB
** negPSRR: 47 dB
** posPSRR: 156 dB
** VoutMax: 3.92001 V
** VoutMin: 0.320001 V
** VcmMax: 3.83001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -8.37529e+07 muA
** NormalTransistorNmos: 4.45581e+07 muA
** NormalTransistorNmos: 4.45571e+07 muA
** NormalTransistorNmos: 4.45581e+07 muA
** NormalTransistorNmos: 4.45571e+07 muA
** NormalTransistorPmos: -8.91179e+07 muA
** NormalTransistorPmos: -4.45589e+07 muA
** NormalTransistorPmos: -4.45589e+07 muA
** NormalTransistorNmos: 1.10227e+08 muA
** NormalTransistorNmos: 1.10226e+08 muA
** NormalTransistorPmos: -1.10226e+08 muA
** NormalTransistorPmos: -1.10227e+08 muA
** DiodeTransistorPmos: -1.092e+08 muA
** DiodeTransistorPmos: -1.09201e+08 muA
** NormalTransistorNmos: 1.09201e+08 muA
** NormalTransistorNmos: 1.092e+08 muA
** DiodeTransistorNmos: 8.37521e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17901  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 4.09501  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 2.78201  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.721001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.41001  V
** innerStageBias: 3.52001  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END