** Name: two_stage_single_output_op_amp_48_7

.MACRO two_stage_single_output_op_amp_48_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=9e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=84e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=18e-6
m4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
m5 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=598e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=598e-6
m7 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=150e-6
m8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=150e-6
m9 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=160e-6
m10 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=160e-6
m11 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=354e-6
m12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=598e-6
m13 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=105e-6
m14 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=384e-6
m15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=294e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=294e-6
m18 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=600e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 19e-12
.EOM two_stage_single_output_op_amp_48_7

** Expected Performance Values: 
** Gain: 111 dB
** Power consumption: 13.4221 mW
** Area: 14524 (mu_m)^2
** Transit frequency: 5.20401 MHz
** Transit frequency with error factor: 5.20344 MHz
** Slew rate: 12.6398 V/mu_s
** Phase margin: 60.1606°
** CMRR: 130 dB
** VoutMax: 4.5 V
** VoutMin: 0.170001 V
** VcmMax: 3.59001 V
** VcmMin: -0.389999 V


** Expected Currents: 
** NormalTransistorPmos: -5.91559e+07 muA
** NormalTransistorPmos: -2.15607e+08 muA
** NormalTransistorNmos: 2.42868e+08 muA
** NormalTransistorNmos: 4.11885e+08 muA
** NormalTransistorNmos: 2.42869e+08 muA
** NormalTransistorNmos: 4.11886e+08 muA
** DiodeTransistorPmos: -2.42867e+08 muA
** NormalTransistorPmos: -2.42868e+08 muA
** NormalTransistorPmos: -2.42868e+08 muA
** DiodeTransistorPmos: -2.42868e+08 muA
** NormalTransistorPmos: -3.38034e+08 muA
** NormalTransistorPmos: -1.69017e+08 muA
** NormalTransistorPmos: -1.69017e+08 muA
** NormalTransistorNmos: 1.56592e+09 muA
** NormalTransistorPmos: -1.56591e+09 muA
** DiodeTransistorNmos: 5.91551e+07 muA
** DiodeTransistorNmos: 2.15608e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.93601  V
** outVoltageBiasXXnXX1: 1.14501  V
** outVoltageBiasXXnXX2: 0.580001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.28601  V
** innerTransistorStack1Load2: 4.28601  V
** out1: 3.57201  V
** sourceGCC1: 0.375  V
** sourceGCC2: 0.375  V
** sourceTransconductance: 3.60001  V


.END