** Name: two_stage_single_output_op_amp_64_2

.MACRO two_stage_single_output_op_amp_64_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=98e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=12e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=29e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=573e-6
m6 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=446e-6
m7 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=135e-6
m8 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=600e-6
m9 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=464e-6
m10 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=16e-6
m11 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=464e-6
m12 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=467e-6
m13 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=467e-6
m14 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=517e-6
m15 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=112e-6
m16 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=582e-6
m17 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=446e-6
m18 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=67e-6
m19 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=135e-6
m20 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=61e-6
m21 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=61e-6
m22 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=573e-6
m23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=29e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 14.4001e-12
.EOM two_stage_single_output_op_amp_64_2

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 7.86401 mW
** Area: 14991 (mu_m)^2
** Transit frequency: 6.25801 MHz
** Transit frequency with error factor: 6.25776 MHz
** Slew rate: 14.2114 V/mu_s
** Phase margin: 60.1606°
** CMRR: 129 dB
** VoutMax: 4.63001 V
** VoutMin: 0.320001 V
** VcmMax: 3 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.52381e+07 muA
** NormalTransistorPmos: -5.66889e+07 muA
** NormalTransistorPmos: -9.33279e+07 muA
** NormalTransistorNmos: 2.94584e+08 muA
** NormalTransistorNmos: 4.47546e+08 muA
** NormalTransistorNmos: 2.94584e+08 muA
** NormalTransistorNmos: 4.47546e+08 muA
** DiodeTransistorPmos: -2.94583e+08 muA
** DiodeTransistorPmos: -2.94584e+08 muA
** NormalTransistorPmos: -2.94583e+08 muA
** NormalTransistorPmos: -2.94584e+08 muA
** NormalTransistorPmos: -3.05926e+08 muA
** DiodeTransistorPmos: -3.05927e+08 muA
** NormalTransistorPmos: -1.52962e+08 muA
** NormalTransistorPmos: -1.52962e+08 muA
** NormalTransistorNmos: 4.92442e+08 muA
** NormalTransistorNmos: 4.92441e+08 muA
** NormalTransistorPmos: -4.92439e+08 muA
** DiodeTransistorNmos: 5.66881e+07 muA
** DiodeTransistorNmos: 9.33271e+07 muA
** DiodeTransistorPmos: -1.52389e+07 muA
** NormalTransistorPmos: -1.52399e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.06101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.52801  V
** outSourceVoltageBiasXXpXX1: 4.26401  V
** outVoltageBiasXXnXX1: 0.905001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 2.93001  V
** innerTransistorStack1Load2: 3.82801  V
** innerTransistorStack2Load2: 3.82601  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.59201  V
** innerTransconductance: 0.329001  V
** inner: 4.26301  V


.END