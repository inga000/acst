.suckt  two_stage_fully_differential_op_amp_27_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_3 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_4 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_5 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_Load_6 outFeedback outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_8 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackStage_Transconductor_9 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_11 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FeedbackStage_Transconductor_12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FirstStage_Load_13 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_14 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_StageBias_15 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_FullyDifferential_FirstStage_StageBias_16 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Transconductor_17 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_FullyDifferential_FirstStage_Transconductor_18 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_Transconductor_19 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m_FullyDifferential_SecondStage1_Transconductor_20 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_21 out1 outVoltageBiasXXpXX2 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m_FullyDifferential_SecondStage1_StageBias_22 SecondStage1YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_Transconductor_23 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m_FullyDifferential_SecondStage2_Transconductor_24 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_StageBias_25 out2 outVoltageBiasXXpXX2 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m_FullyDifferential_SecondStage2_StageBias_26 SecondStage2YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_27 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_28 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_29 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_FullyDifferential_MainBias_30 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_31 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_32 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_27_4

