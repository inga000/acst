** Name: symmetrical_op_amp147

.MACRO symmetrical_op_amp147 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=31e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias3 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=112e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=6e-6 W=112e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=251e-6
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=251e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=272e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=272e-6
mSymmetricalFirstStageLoad10 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=61e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=1e-6 W=24e-6
mSecondStage1Transconductor12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=24e-6
mSymmetricalFirstStageLoad13 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=61e-6
mSymmetricalFirstStageStageBias14 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=315e-6
mSymmetricalFirstStageStageBias15 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=158e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias16 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=112e-6
mSymmetricalFirstStageTransconductor17 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=238e-6
mSecondStage1StageBias18 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=6e-6 W=112e-6
mSymmetricalFirstStageTransconductor19 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=238e-6
mMainBias20 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=506e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp147

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 5.99901 mW
** Area: 7502 (mu_m)^2
** Transit frequency: 14.1901 MHz
** Transit frequency with error factor: 14.1904 MHz
** Slew rate: 17.342 V/mu_s
** Phase margin: 70.4739°
** CMRR: 142 dB
** negPSRR: 47 dB
** posPSRR: 53 dB
** VoutMax: 3 V
** VoutMin: 0.440001 V
** VcmMax: 3.11001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -5.13021e+08 muA
** NormalTransistorNmos: 1.59686e+08 muA
** NormalTransistorNmos: 1.59685e+08 muA
** NormalTransistorNmos: 1.59686e+08 muA
** NormalTransistorNmos: 1.59685e+08 muA
** NormalTransistorPmos: -3.19371e+08 muA
** NormalTransistorPmos: -3.1937e+08 muA
** NormalTransistorPmos: -1.59685e+08 muA
** NormalTransistorPmos: -1.59685e+08 muA
** NormalTransistorNmos: 1.73702e+08 muA
** NormalTransistorNmos: 1.73701e+08 muA
** NormalTransistorPmos: -1.73701e+08 muA
** DiodeTransistorPmos: -1.73701e+08 muA
** DiodeTransistorPmos: -1.73702e+08 muA
** NormalTransistorPmos: -1.73701e+08 muA
** NormalTransistorNmos: 1.73703e+08 muA
** NormalTransistorNmos: 1.73702e+08 muA
** DiodeTransistorNmos: 5.13022e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 3.71801  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 2.43601  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.846001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.29701  V
** innerTransistorStack1Load1: 0.265001  V
** innerTransistorStack2Load1: 0.265001  V
** sourceTransconductance: 3.25701  V
** innerTransconductance: 0.150001  V
** inner: 3.71901  V
** inner: 0.150001  V


.END