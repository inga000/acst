.suckt  two_stage_single_output_op_amp_3_5 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m4 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
m5 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m6 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourceNmos sourceNmos nmos
m7 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c2 out sourceNmos 
m10 out outFirstStage sourceNmos sourceNmos nmos
m11 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m12 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m13 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m14 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m15 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m17 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_3_5

