** Name: one_stage_single_output_op_amp65

.MACRO one_stage_single_output_op_amp65 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=10e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
m3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
m4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
m5 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=145e-6
m6 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=45e-6
m7 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
m8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=145e-6
m9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=433e-6
m10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=433e-6
m11 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=190e-6
m12 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=292e-6
m13 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=257e-6
m14 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=257e-6
m15 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=190e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=346e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=346e-6
m18 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=173e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp65

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 3.08401 mW
** Area: 7742 (mu_m)^2
** Transit frequency: 7.05001 MHz
** Transit frequency with error factor: 7.05046 MHz
** Slew rate: 9.32819 V/mu_s
** Phase margin: 87.0896°
** CMRR: 139 dB
** VoutMax: 4.47001 V
** VoutMin: 0.770001 V
** VcmMax: 3.11001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.00231e+07 muA
** NormalTransistorNmos: 1.04641e+07 muA
** NormalTransistorNmos: 1.87255e+08 muA
** NormalTransistorNmos: 2.83177e+08 muA
** NormalTransistorNmos: 1.87255e+08 muA
** NormalTransistorNmos: 2.83177e+08 muA
** NormalTransistorPmos: -1.87254e+08 muA
** NormalTransistorPmos: -1.87255e+08 muA
** NormalTransistorPmos: -1.87254e+08 muA
** NormalTransistorPmos: -1.87255e+08 muA
** NormalTransistorPmos: -1.91846e+08 muA
** NormalTransistorPmos: -1.91847e+08 muA
** NormalTransistorPmos: -9.59229e+07 muA
** NormalTransistorPmos: -9.59229e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.00239e+07 muA
** DiodeTransistorPmos: -1.04649e+07 muA


** Expected Voltages: 
** ibias: 1.15101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.24401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.60101  V
** innerTransistorStack1Load2: 4.58101  V
** innerTransistorStack2Load2: 4.58101  V
** out1: 4.23401  V
** sourceGCC1: 0.531001  V
** sourceGCC2: 0.531001  V
** sourceTransconductance: 3.27901  V


.END