.suckt  symmetrical_op_amp191 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m2 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m3 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m4 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m5 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
m6 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m8 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m9 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m10 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m11 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m12 out outVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m13 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
m14 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m16 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
m17 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m19 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m20 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m21 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m22 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m23 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos
.end symmetrical_op_amp191

