.suckt  two_stage_fully_differential_op_amp_67_6 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m3 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m4 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m5 inputVoltageBiasXXnXX4 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m6 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m7 outFeedback outFeedback sourcePmos sourcePmos pmos
m8 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m9 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m14 out1FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m15 out2FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m16 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m17 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m18 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m19 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m20 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m21 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m22 out1 outVoltageBiasXXnXX3 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m23 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m24 out1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m25 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m26 out2 outVoltageBiasXXnXX3 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m27 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m28 out2 ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m29 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m30 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m31 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m32 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos
m33 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m34 inputVoltageBiasXXnXX4 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m35 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m36 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m37 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m38 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_67_6

