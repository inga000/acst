** Name: two_stage_single_output_op_amp_47_5

.MACRO two_stage_single_output_op_amp_47_5 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=13e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
m3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=74e-6
m4 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=9e-6 W=147e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=23e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=484e-6
m7 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=391e-6
m8 inputVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=22e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=63e-6
m10 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=20e-6
m11 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=105e-6
m12 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=20e-6
m13 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=77e-6
m14 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=77e-6
m15 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=484e-6
m16 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=202e-6
m17 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=202e-6
m18 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=29e-6
m19 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=29e-6
m20 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=15e-6
m21 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=15e-6
m22 FirstStageYsourceTransconductance inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=9e-6 W=350e-6
m23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_47_5

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 5.52101 mW
** Area: 12020 (mu_m)^2
** Transit frequency: 3.60301 MHz
** Transit frequency with error factor: 3.60272 MHz
** Slew rate: 4.28673 V/mu_s
** Phase margin: 71.0468°
** CMRR: 135 dB
** VoutMax: 3.81001 V
** VoutMin: 0.560001 V
** VcmMax: 4.08001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.99981e+07 muA
** NormalTransistorNmos: 1.5027e+08 muA
** NormalTransistorNmos: 8.38101e+06 muA
** NormalTransistorNmos: 1.94721e+07 muA
** NormalTransistorNmos: 2.93321e+07 muA
** NormalTransistorNmos: 1.94721e+07 muA
** NormalTransistorNmos: 2.93321e+07 muA
** NormalTransistorPmos: -1.94729e+07 muA
** NormalTransistorPmos: -1.94739e+07 muA
** NormalTransistorPmos: -1.94729e+07 muA
** NormalTransistorPmos: -1.94739e+07 muA
** NormalTransistorPmos: -1.97229e+07 muA
** NormalTransistorPmos: -9.86099e+06 muA
** NormalTransistorPmos: -9.86099e+06 muA
** NormalTransistorNmos: 8.36823e+08 muA
** NormalTransistorPmos: -8.36822e+08 muA
** DiodeTransistorPmos: -8.36823e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.99989e+07 muA
** NormalTransistorPmos: -4e+07 muA
** DiodeTransistorPmos: -1.50269e+08 muA
** DiodeTransistorPmos: -8.38199e+06 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.68601  V
** inputVoltageBiasXXpXX3: 4.26701  V
** out: 2.5  V
** outFirstStage: 0.968001  V
** outInputVoltageBiasXXpXX1: 3.24801  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.12401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.05001  V
** innerTransistorStack1Load2: 4.41401  V
** innerTransistorStack2Load2: 4.41401  V
** sourceGCC1: 0.527001  V
** sourceGCC2: 0.527001  V
** sourceTransconductance: 3.25501  V
** inner: 4.12301  V


.END