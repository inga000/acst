.suckt  two_stage_single_output_op_amp_37_4 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m4 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m5 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos
m6 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m7 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos
m8 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m9 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c2 out sourceNmos 
m12 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m13 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m14 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m15 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m16 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m17 ibias ibias sourceNmos sourceNmos nmos
m18 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m19 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_37_4

