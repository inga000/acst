** Name: symmetrical_op_amp115

.MACRO symmetrical_op_amp115 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=1e-6 W=18e-6
mMainBias4 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=66e-6
mSecondStage1StageBias6 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mSymmetricalFirstStageTransconductor7 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=35e-6
mSecondStage1StageBias8 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=21e-6
mSymmetricalFirstStageTransconductor9 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=35e-6
mMainBias10 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=3e-6 W=99e-6
mSymmetricalFirstStageLoad11 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=46e-6
mSymmetricalFirstStageLoad12 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=46e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=57e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=57e-6
mSymmetricalFirstStageLoad15 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=81e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=102e-6
mSecondStage1Transconductor17 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=102e-6
mSymmetricalFirstStageLoad18 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=81e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp115

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 1.28501 mW
** Area: 3176 (mu_m)^2
** Transit frequency: 2.73701 MHz
** Transit frequency with error factor: 2.73671 MHz
** Slew rate: 4.11001 V/mu_s
** Phase margin: 80.2142°
** CMRR: 141 dB
** negPSRR: 120 dB
** posPSRR: 61 dB
** VoutMax: 4.25 V
** VoutMin: 0.730001 V
** VcmMax: 4.81001 V
** VcmMin: 0.830001 V


** Expected Currents: 
** NormalTransistorNmos: 9.96151e+07 muA
** NormalTransistorPmos: -3.25859e+07 muA
** NormalTransistorPmos: -3.25869e+07 muA
** NormalTransistorPmos: -3.25859e+07 muA
** NormalTransistorPmos: -3.25869e+07 muA
** NormalTransistorNmos: 6.51701e+07 muA
** NormalTransistorNmos: 3.25851e+07 muA
** NormalTransistorNmos: 3.25851e+07 muA
** NormalTransistorNmos: 4.11551e+07 muA
** NormalTransistorNmos: 4.11541e+07 muA
** NormalTransistorPmos: -4.11559e+07 muA
** NormalTransistorPmos: -4.11549e+07 muA
** DiodeTransistorNmos: 4.11531e+07 muA
** DiodeTransistorNmos: 4.11521e+07 muA
** NormalTransistorPmos: -4.11539e+07 muA
** NormalTransistorPmos: -4.11549e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.96159e+07 muA


** Expected Voltages: 
** ibias: 0.593001  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 0.579001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 1.14801  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.86001  V
** innerStageBias: 0.591001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END