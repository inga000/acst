** Name: two_stage_single_output_op_amp_63_2

.MACRO two_stage_single_output_op_amp_63_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=57e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=57e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mMainBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=141e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=509e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=509e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=532e-6
mMainBias11 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=407e-6
mSecondStage1Transconductor12 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=532e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=141e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=320e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=57e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=332e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=332e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=600e-6
mMainBias19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=70e-6
mSecondStage1StageBias20 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=57e-6
mMainBias22 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14e-12
.EOM two_stage_single_output_op_amp_63_2

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 7.51001 mW
** Area: 14998 (mu_m)^2
** Transit frequency: 7.64201 MHz
** Transit frequency with error factor: 7.6421 MHz
** Slew rate: 13.4005 V/mu_s
** Phase margin: 60.1606°
** CMRR: 119 dB
** VoutMax: 4.69001 V
** VoutMin: 0.300001 V
** VcmMax: 3.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.61005e+08 muA
** NormalTransistorPmos: -5.91559e+07 muA
** NormalTransistorPmos: -8.28399e+06 muA
** NormalTransistorNmos: 1.88593e+08 muA
** NormalTransistorNmos: 3.23303e+08 muA
** NormalTransistorNmos: 1.88589e+08 muA
** NormalTransistorNmos: 3.23297e+08 muA
** DiodeTransistorPmos: -1.8859e+08 muA
** DiodeTransistorPmos: -1.88589e+08 muA
** NormalTransistorPmos: -1.88588e+08 muA
** NormalTransistorPmos: -1.88589e+08 muA
** NormalTransistorPmos: -2.69418e+08 muA
** NormalTransistorPmos: -2.69419e+08 muA
** NormalTransistorPmos: -1.34708e+08 muA
** NormalTransistorPmos: -1.34708e+08 muA
** NormalTransistorNmos: 5.07054e+08 muA
** NormalTransistorNmos: 5.07053e+08 muA
** NormalTransistorPmos: -5.07052e+08 muA
** DiodeTransistorNmos: 5.91551e+07 muA
** DiodeTransistorNmos: 8.28301e+06 muA
** DiodeTransistorPmos: -2.61004e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.932001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40801  V
** innerTransistorStack1Load2: 3.68801  V
** innerTransistorStack2Load2: 3.68101  V
** out1: 2.375  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.46101  V
** innerTransconductance: 0.377001  V


.END