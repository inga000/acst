** Name: two_stage_single_output_op_amp_8_12

.MACRO two_stage_single_output_op_amp_8_12 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=19e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=33e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=72e-6
m4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=13e-6
m5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=315e-6
m7 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=72e-6
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=195e-6
m9 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=46e-6
m10 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=194e-6
m11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=195e-6
m12 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=324e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=33e-6
m14 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
m15 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=315e-6
m16 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=358e-6
m17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=543e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 11.5e-12
.EOM two_stage_single_output_op_amp_8_12

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 11.9141 mW
** Area: 14940 (mu_m)^2
** Transit frequency: 10.7251 MHz
** Transit frequency with error factor: 10.7074 MHz
** Slew rate: 14.3925 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** negPSRR: 165 dB
** posPSRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 1.77001 V
** VcmMax: 4.47001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorNmos: 2.38571e+07 muA
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -6.45106e+08 muA
** DiodeTransistorPmos: -8.36689e+07 muA
** NormalTransistorPmos: -8.36689e+07 muA
** NormalTransistorNmos: 1.67338e+08 muA
** NormalTransistorNmos: 8.36681e+07 muA
** NormalTransistorNmos: 8.36681e+07 muA
** NormalTransistorNmos: 1.43498e+09 muA
** DiodeTransistorNmos: 1.43497e+09 muA
** NormalTransistorPmos: -1.43497e+09 muA
** NormalTransistorPmos: -1.43497e+09 muA
** DiodeTransistorNmos: 6.45107e+08 muA
** NormalTransistorNmos: 6.45107e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.38579e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 0.562001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.05001  V
** outInputVoltageBiasXXnXX1: 2.17601  V
** outSourceVoltageBiasXXnXX1: 1.08801  V
** outVoltageBiasXXpXX0: 3.72301  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.06901  V
** sourceTransconductance: 1.88101  V
** innerTransconductance: 4.61401  V
** inner: 1.08801  V


.END