** Name: two_stage_single_output_op_amp_55_1

.MACRO two_stage_single_output_op_amp_55_1 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=20e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=20e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=10e-6 W=50e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=31e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=54e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=20e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=20e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=20e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=10e-6 W=105e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=69e-6
mFoldedCascodeFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=8e-6 W=20e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=529e-6
mMainBias13 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=288e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=35e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mSecondStage1StageBias17 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=573e-6
mFoldedCascodeFirstStageLoad18 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=35e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_55_1

** Expected Performance Values: 
** Gain: 115 dB
** Power consumption: 4.20101 mW
** Area: 11662 (mu_m)^2
** Transit frequency: 3.52001 MHz
** Transit frequency with error factor: 3.51986 MHz
** Slew rate: 4.21999 V/mu_s
** Phase margin: 61.8795°
** CMRR: 134 dB
** VoutMax: 4.76001 V
** VoutMin: 0.650001 V
** VcmMax: 5.16001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorNmos: 1.04918e+08 muA
** NormalTransistorNmos: 5.75551e+07 muA
** NormalTransistorPmos: -1.90469e+07 muA
** NormalTransistorPmos: -2.93479e+07 muA
** NormalTransistorPmos: -1.90469e+07 muA
** NormalTransistorPmos: -2.93479e+07 muA
** DiodeTransistorNmos: 1.90461e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90461e+07 muA
** DiodeTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 2.06011e+07 muA
** NormalTransistorNmos: 1.03001e+07 muA
** NormalTransistorNmos: 1.03001e+07 muA
** NormalTransistorNmos: 6.08955e+08 muA
** NormalTransistorPmos: -6.08954e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.04917e+08 muA
** DiodeTransistorPmos: -5.75559e+07 muA


** Expected Voltages: 
** ibias: 0.558001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 1.05401  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.19301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.553001  V
** out1: 1.25901  V
** sourceGCC1: 4.55101  V
** sourceGCC2: 4.55101  V
** sourceTransconductance: 1.88801  V


.END