** Name: two_stage_single_output_op_amp_75_10

.MACRO two_stage_single_output_op_amp_75_10 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=18e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=14e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=15e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=97e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=24e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=6e-6 W=18e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=18e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=18e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=45e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=377e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=17e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=185e-6
mMainBias14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=31e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=108e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=108e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=197e-6
mMainBias19 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=521e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=410e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=39e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_75_10

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 2.98301 mW
** Area: 5004 (mu_m)^2
** Transit frequency: 4.02801 MHz
** Transit frequency with error factor: 4.0276 MHz
** Slew rate: 3.50745 V/mu_s
** Phase margin: 62.4525°
** CMRR: 144 dB
** VoutMax: 4.53001 V
** VoutMin: 0.160001 V
** VcmMax: 5.25 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 1.31994e+08 muA
** NormalTransistorNmos: 2.21311e+07 muA
** NormalTransistorPmos: -1.17292e+08 muA
** NormalTransistorPmos: -1.58389e+07 muA
** NormalTransistorPmos: -2.44109e+07 muA
** NormalTransistorPmos: -1.58389e+07 muA
** NormalTransistorPmos: -2.44109e+07 muA
** DiodeTransistorNmos: 1.58381e+07 muA
** NormalTransistorNmos: 1.58381e+07 muA
** NormalTransistorNmos: 1.58381e+07 muA
** NormalTransistorNmos: 1.71421e+07 muA
** NormalTransistorNmos: 1.71411e+07 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 8.57101e+06 muA
** NormalTransistorNmos: 2.6627e+08 muA
** NormalTransistorPmos: -2.66269e+08 muA
** NormalTransistorPmos: -2.6627e+08 muA
** DiodeTransistorNmos: 1.17293e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.31993e+08 muA
** DiodeTransistorPmos: -2.21319e+07 muA


** Expected Voltages: 
** ibias: 0.564001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.08801  V
** out: 2.5  V
** outFirstStage: 4.16001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.27701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.533001  V
** innerTransistorStack2Load2: 0.449001  V
** out1: 0.654001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.44001  V


.END