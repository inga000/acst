.suckt  two_stage_single_output_op_amp_149_4 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m4 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m5 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos
m6 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos
m8 FirstStageYinnerSourceLoad1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m9 outFirstStage outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m11 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c2 out sourceNmos 
m13 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m14 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m15 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m16 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m17 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m18 ibias ibias sourceNmos sourceNmos nmos
m19 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m20 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_149_4

