.suckt  two_stage_fully_differential_op_amp_69_7 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m3 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m4 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m5 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m6 outFeedback outFeedback sourcePmos sourcePmos pmos
m7 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m8 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m9 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m14 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m15 out1FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m16 FirstStageYinnerTransistorStack1Load2 outFeedback sourcePmos sourcePmos pmos
m17 out2FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m18 FirstStageYinnerTransistorStack2Load2 outFeedback sourcePmos sourcePmos pmos
m19 sourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m20 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m21 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m22 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m23 out1 ibias sourceNmos sourceNmos nmos
m24 out1 out1FirstStage sourcePmos sourcePmos pmos
m25 out2 ibias sourceNmos sourceNmos nmos
m26 out2 out2FirstStage sourcePmos sourcePmos pmos
m27 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
m28 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m29 ibias ibias sourceNmos sourceNmos nmos
m30 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m31 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_69_7

