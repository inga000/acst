** Name: two_stage_single_output_op_amp_24_5

.MACRO two_stage_single_output_op_amp_24_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=160e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=61e-6
mMainBias3 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=3e-6 W=20e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=281e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=124e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=414e-6
mSimpleFirstStageLoad7 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=5e-6 W=132e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=105e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=105e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=443e-6
mSimpleFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=132e-6
mMainBias12 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=296e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=22e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=124e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=281e-6
mMainBias16 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mMainBias17 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=477e-6
mSecondStage1StageBias18 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=3e-6 W=414e-6
mSimpleFirstStageTransconductor19 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=22e-6
mMainBias20 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=93e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_24_5

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 4.24001 mW
** Area: 11685 (mu_m)^2
** Transit frequency: 4.88801 MHz
** Transit frequency with error factor: 4.87966 MHz
** Slew rate: 7.20203 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 101 dB
** posPSRR: 210 dB
** VoutMax: 3.85001 V
** VoutMin: 0.150001 V
** VcmMax: 3.09001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.27686e+08 muA
** NormalTransistorPmos: -4.73839e+07 muA
** NormalTransistorPmos: -2.41379e+08 muA
** NormalTransistorNmos: 5.02851e+07 muA
** NormalTransistorNmos: 5.02841e+07 muA
** NormalTransistorNmos: 5.02831e+07 muA
** NormalTransistorNmos: 5.02841e+07 muA
** NormalTransistorPmos: -1.00566e+08 muA
** DiodeTransistorPmos: -1.00567e+08 muA
** NormalTransistorPmos: -5.02839e+07 muA
** NormalTransistorPmos: -5.02839e+07 muA
** NormalTransistorNmos: 2.10939e+08 muA
** NormalTransistorPmos: -2.10937e+08 muA
** DiodeTransistorPmos: -2.10936e+08 muA
** DiodeTransistorNmos: 4.73831e+07 muA
** DiodeTransistorNmos: 2.4138e+08 muA
** DiodeTransistorPmos: -2.27685e+08 muA
** NormalTransistorPmos: -2.27686e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.28801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.44401  V
** outSourceVoltageBiasXXpXX1: 4.22201  V
** outSourceVoltageBiasXXpXX2: 4.14501  V
** outVoltageBiasXXnXX0: 0.619001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.42001  V
** inner: 4.22001  V
** inner: 4.14101  V


.END