** Name: two_stage_single_output_op_amp_43_11

.MACRO two_stage_single_output_op_amp_43_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=10e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=179e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=94e-6
mSecondStage1StageBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=67e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=34e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=66e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=66e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=586e-6
mMainBias10 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=324e-6
mSecondStage1StageBias11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=295e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=34e-6
mMainBias13 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=173e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=389e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=600e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=179e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.5e-12
.EOM two_stage_single_output_op_amp_43_11

** Expected Performance Values: 
** Gain: 135 dB
** Power consumption: 6.02801 mW
** Area: 8588 (mu_m)^2
** Transit frequency: 4.625 MHz
** Transit frequency with error factor: 4.61986 MHz
** Slew rate: 5.04307 V/mu_s
** Phase margin: 60.1606°
** CMRR: 100 dB
** VoutMax: 4.25 V
** VoutMin: 0.770001 V
** VcmMax: 3.83001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.70069e+08 muA
** NormalTransistorNmos: 3.18121e+08 muA
** NormalTransistorNmos: 4.31381e+07 muA
** NormalTransistorNmos: 6.47451e+07 muA
** NormalTransistorNmos: 4.31381e+07 muA
** NormalTransistorNmos: 6.47451e+07 muA
** DiodeTransistorPmos: -4.31389e+07 muA
** NormalTransistorPmos: -4.31389e+07 muA
** NormalTransistorPmos: -4.32169e+07 muA
** NormalTransistorPmos: -2.16079e+07 muA
** NormalTransistorPmos: -2.16079e+07 muA
** NormalTransistorNmos: 5.77915e+08 muA
** NormalTransistorNmos: 5.77914e+08 muA
** NormalTransistorPmos: -5.77914e+08 muA
** NormalTransistorPmos: -5.77915e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.70068e+08 muA
** DiodeTransistorPmos: -3.1812e+08 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.00301  V
** out: 2.5  V
** outFirstStage: 4.14801  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.15101  V
** sourceGCC1: 0.537001  V
** sourceGCC2: 0.537001  V
** sourceTransconductance: 3.23701  V
** innerStageBias: 0.495001  V
** innerTransconductance: 4.71201  V


.END