** Name: symmetrical_op_amp14

.MACRO symmetrical_op_amp14 ibias in1 in2 out sourceNmos sourcePmos
m1 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
m2 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
m3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
m5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=75e-6
m6 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=1e-6 W=75e-6
m7 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=13e-6
m8 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=13e-6
m9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=54e-6
m10 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=54e-6
m11 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=25e-6
m12 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=4e-6 W=196e-6
m13 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=75e-6
m14 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=25e-6
m15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=106e-6
m16 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=75e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp14

** Expected Performance Values: 
** Gain: 95 dB
** Power consumption: 0.840001 mW
** Area: 2810 (mu_m)^2
** Transit frequency: 3.32601 MHz
** Transit frequency with error factor: 3.32572 MHz
** Slew rate: 3.58136 V/mu_s
** Phase margin: 69.9009°
** CMRR: 145 dB
** negPSRR: 48 dB
** posPSRR: 52 dB
** VoutMax: 4.11001 V
** VoutMin: 0.660001 V
** VcmMax: 4.03001 V
** VcmMin: 0.0600001 V


** Expected Currents: 
** NormalTransistorPmos: -4.93609e+07 muA
** DiodeTransistorNmos: 1.34321e+07 muA
** DiodeTransistorNmos: 1.34321e+07 muA
** NormalTransistorPmos: -2.68669e+07 muA
** NormalTransistorPmos: -1.34329e+07 muA
** NormalTransistorPmos: -1.34329e+07 muA
** NormalTransistorNmos: 3.58471e+07 muA
** NormalTransistorNmos: 3.58481e+07 muA
** NormalTransistorPmos: -3.58479e+07 muA
** DiodeTransistorPmos: -3.58489e+07 muA
** DiodeTransistorPmos: -3.58479e+07 muA
** NormalTransistorPmos: -3.58489e+07 muA
** NormalTransistorNmos: 3.58471e+07 muA
** NormalTransistorNmos: 3.58481e+07 muA
** DiodeTransistorNmos: 4.93601e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 1.06301  V
** inSourceStageBiasComplementarySecondStage: 4.27201  V
** inSourceTransconductanceComplementarySecondStage: 0.623001  V
** innerComplementarySecondStage: 3.54401  V
** out: 2.5  V
** outFirstStage: 0.623001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.23701  V
** innerTransconductance: 0.218001  V
** inner: 4.27101  V
** inner: 0.218001  V


.END