** Name: two_stage_single_output_op_amp_45_5

.MACRO two_stage_single_output_op_amp_45_5 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=11e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=21e-6
m4 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=24e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=9e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=520e-6
m7 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
m8 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=49e-6
m9 inputVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=19e-6
m10 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=22e-6
m11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=36e-6
m12 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=36e-6
m14 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=137e-6
m15 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=137e-6
m16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=520e-6
m17 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=9e-6 W=211e-6
m18 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
m19 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=77e-6
m20 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=77e-6
m21 FirstStageYsourceTransconductance inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=114e-6
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=9e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_45_5

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 3.77501 mW
** Area: 13138 (mu_m)^2
** Transit frequency: 4.03801 MHz
** Transit frequency with error factor: 4.03781 MHz
** Slew rate: 9.55022 V/mu_s
** Phase margin: 63.0254°
** CMRR: 132 dB
** VoutMax: 3.12001 V
** VoutMin: 0.560001 V
** VcmMax: 3.85001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.00001e+07 muA
** NormalTransistorNmos: 2.33321e+07 muA
** NormalTransistorNmos: 9.09201e+06 muA
** NormalTransistorNmos: 4.34491e+07 muA
** NormalTransistorNmos: 6.52341e+07 muA
** NormalTransistorNmos: 4.34491e+07 muA
** NormalTransistorNmos: 6.52341e+07 muA
** DiodeTransistorPmos: -4.34499e+07 muA
** NormalTransistorPmos: -4.34499e+07 muA
** NormalTransistorPmos: -4.34499e+07 muA
** NormalTransistorPmos: -4.35729e+07 muA
** NormalTransistorPmos: -2.17859e+07 muA
** NormalTransistorPmos: -2.17859e+07 muA
** NormalTransistorNmos: 5.72058e+08 muA
** NormalTransistorPmos: -5.72057e+08 muA
** DiodeTransistorPmos: -5.72058e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.00009e+07 muA
** NormalTransistorPmos: -1.00019e+07 muA
** DiodeTransistorPmos: -2.33329e+07 muA
** DiodeTransistorPmos: -9.09299e+06 muA


** Expected Voltages: 
** ibias: 1.16701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.68601  V
** inputVoltageBiasXXpXX3: 4.23001  V
** out: 2.5  V
** outFirstStage: 0.962001  V
** outInputVoltageBiasXXpXX1: 2.55401  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.77701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.57101  V
** out1: 4.20701  V
** sourceGCC1: 0.522001  V
** sourceGCC2: 0.522001  V
** sourceTransconductance: 3.44001  V
** inner: 3.77501  V


.END