.suckt  two_stage_single_output_op_amp_103_6 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_3 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_4 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m_SingleOutput_FirstStage_Load_6 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m_SingleOutput_FirstStage_Load_7 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m_SingleOutput_FirstStage_Load_9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_StageBias_10 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m_SingleOutput_FirstStage_StageBias_11 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Transconductor_12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m_SingleOutput_FirstStage_Transconductor_13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_Transconductor_14 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_SingleOutput_SecondStage1_Transconductor_15 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_SingleOutput_SecondStage1_StageBias_17 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_18 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_19 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_20 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_SingleOutput_MainBias_21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_22 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos
m_SingleOutput_MainBias_23 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos
m_SingleOutput_MainBias_24 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_103_6

