** Name: two_stage_single_output_op_amp_12_7

.MACRO two_stage_single_output_op_amp_12_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mMainBias2 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
mSimpleFirstStageTransconductor3 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=12e-6
mSimpleFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=82e-6
mMainBias5 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=111e-6
mSecondStage1StageBias6 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mSimpleFirstStageTransconductor7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=12e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=28e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=28e-6
mSimpleFirstStageLoad10 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=128e-6
mSecondStage1Transconductor11 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=381e-6
mSimpleFirstStageLoad12 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=128e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_12_7

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 2.37501 mW
** Area: 4582 (mu_m)^2
** Transit frequency: 5.33901 MHz
** Transit frequency with error factor: 5.33621 MHz
** Slew rate: 5.1214 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** negPSRR: 119 dB
** posPSRR: 104 dB
** VoutMax: 4.77001 V
** VoutMin: 0.170001 V
** VcmMax: 5.10001 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 6.43031e+07 muA
** NormalTransistorPmos: -2.36739e+07 muA
** NormalTransistorPmos: -2.36749e+07 muA
** NormalTransistorPmos: -2.36739e+07 muA
** NormalTransistorPmos: -2.36749e+07 muA
** NormalTransistorNmos: 4.73461e+07 muA
** NormalTransistorNmos: 2.36731e+07 muA
** NormalTransistorNmos: 2.36731e+07 muA
** NormalTransistorNmos: 3.53427e+08 muA
** NormalTransistorPmos: -3.53426e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.43039e+07 muA


** Expected Voltages: 
** ibias: 0.571001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.20801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.42601  V
** innerTransistorStack2Load1: 4.42601  V
** out1: 4.12901  V
** sourceTransconductance: 1.94201  V


.END