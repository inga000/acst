** Name: two_stage_single_output_op_amp_55_3

.MACRO two_stage_single_output_op_amp_55_3 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
m2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=24e-6
m3 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=37e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
m6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
m7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=66e-6
m8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=66e-6
m9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=9e-6 W=236e-6
m10 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=400e-6
m11 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=121e-6
m12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=6e-6 W=24e-6
m13 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=68e-6
m14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m16 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=244e-6
m17 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=328e-6
m18 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=68e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 8e-12
.EOM two_stage_single_output_op_amp_55_3

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 10.0221 mW
** Area: 8040 (mu_m)^2
** Transit frequency: 8.31301 MHz
** Transit frequency with error factor: 8.31256 MHz
** Slew rate: 5.69787 V/mu_s
** Phase margin: 60.1606°
** CMRR: 137 dB
** VoutMax: 3.27001 V
** VoutMin: 0.720001 V
** VcmMax: 4.78001 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorNmos: 1.07123e+08 muA
** NormalTransistorPmos: -4.57119e+07 muA
** NormalTransistorPmos: -7.71399e+07 muA
** NormalTransistorPmos: -4.57119e+07 muA
** NormalTransistorPmos: -7.71399e+07 muA
** DiodeTransistorNmos: 4.57111e+07 muA
** NormalTransistorNmos: 4.57121e+07 muA
** NormalTransistorNmos: 4.57111e+07 muA
** DiodeTransistorNmos: 4.57121e+07 muA
** NormalTransistorNmos: 6.28531e+07 muA
** NormalTransistorNmos: 3.14271e+07 muA
** NormalTransistorNmos: 3.14271e+07 muA
** NormalTransistorNmos: 1.73299e+09 muA
** NormalTransistorPmos: -1.73298e+09 muA
** NormalTransistorPmos: -1.73299e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.07122e+08 muA
** DiodeTransistorPmos: -1.07121e+08 muA


** Expected Voltages: 
** ibias: 0.574001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 2.50201  V
** out: 2.5  V
** outFirstStage: 1.12101  V
** outSourceVoltageBiasXXpXX1: 3.80701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.552001  V
** out1: 1.32601  V
** sourceGCC1: 3.25901  V
** sourceGCC2: 3.25901  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 3.60801  V


.END