** Name: two_stage_single_output_op_amp_114_10

.MACRO two_stage_single_output_op_amp_114_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=11e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=20e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=413e-6
m4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=494e-6
m5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
m6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
m7 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=279e-6
m8 out ibias sourceNmos sourceNmos nmos4 L=7e-6 W=349e-6
m9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=16e-6
m10 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=47e-6
m11 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=45e-6
m12 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=413e-6
m13 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=47e-6
m14 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=66e-6
m15 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=7e-6 W=66e-6
m16 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
m17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=549e-6
m18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=279e-6
m19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=13e-6
m20 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=259e-6
m21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=546e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10.4001e-12
.EOM two_stage_single_output_op_amp_114_10

** Expected Performance Values: 
** Gain: 107 dB
** Power consumption: 6.00601 mW
** Area: 14903 (mu_m)^2
** Transit frequency: 3.63401 MHz
** Transit frequency with error factor: 3.63212 MHz
** Slew rate: 10.1792 V/mu_s
** Phase margin: 60.1606°
** CMRR: 80 dB
** VoutMax: 4.57001 V
** VoutMin: 0.270001 V
** VcmMax: 4.52001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 1.45651e+07 muA
** NormalTransistorNmos: 4.01561e+07 muA
** NormalTransistorPmos: -3.83939e+07 muA
** NormalTransistorPmos: -7.50694e+08 muA
** NormalTransistorNmos: 1.79571e+07 muA
** NormalTransistorNmos: 1.79571e+07 muA
** DiodeTransistorPmos: -1.79579e+07 muA
** NormalTransistorPmos: -1.79579e+07 muA
** NormalTransistorNmos: 7.86612e+08 muA
** DiodeTransistorNmos: 7.86612e+08 muA
** NormalTransistorNmos: 1.79581e+07 muA
** NormalTransistorNmos: 1.79581e+07 muA
** NormalTransistorNmos: 3.1143e+08 muA
** NormalTransistorPmos: -3.11429e+08 muA
** NormalTransistorPmos: -3.1143e+08 muA
** DiodeTransistorNmos: 3.83931e+07 muA
** NormalTransistorNmos: 3.83921e+07 muA
** DiodeTransistorNmos: 7.50695e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.45659e+07 muA
** DiodeTransistorPmos: -4.01569e+07 muA


** Expected Voltages: 
** ibias: 0.678001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.62701  V
** out: 2.5  V
** outFirstStage: 4.25701  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX1: 3.48401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.26601  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 4.29901  V
** inner: 0.554001  V


.END