.suckt  one_stage_fully_differential_op_amp50 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
m1 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m2 outFeedback outFeedback sourcePmos sourcePmos pmos
m3 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m4 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m5 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m6 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m7 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m8 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m9 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m10 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m11 out1 outFeedback sourcePmos sourcePmos pmos
m12 out2 outFeedback sourcePmos sourcePmos pmos
m13 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m14 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m15 out1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m16 out2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out1 sourceNmos 
c2 out2 sourceNmos 
m17 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m18 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
.end one_stage_fully_differential_op_amp50

