** Name: two_stage_single_output_op_amp_106_1

.MACRO two_stage_single_output_op_amp_106_1 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=34e-6
m2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=10e-6 W=71e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=10e-6 W=71e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=24e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=39e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=346e-6
m7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=6e-6
m8 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=182e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=71e-6
m10 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=11e-6
m11 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=41e-6
m12 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=10e-6 W=71e-6
m13 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=40e-6
m14 out ibias sourcePmos sourcePmos pmos4 L=6e-6 W=543e-6
m15 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=5e-6 W=9e-6
m16 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=346e-6
m17 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=5e-6 W=9e-6
m18 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=81e-6
m19 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=81e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=39e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.30001e-12
.EOM two_stage_single_output_op_amp_106_1

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 1.59701 mW
** Area: 14992 (mu_m)^2
** Transit frequency: 2.65701 MHz
** Transit frequency with error factor: 2.65717 MHz
** Slew rate: 7.49447 V/mu_s
** Phase margin: 60.1606°
** CMRR: 136 dB
** VoutMax: 4.63001 V
** VoutMin: 0.300001 V
** VcmMax: 3.15001 V
** VcmMin: 1.20001 V


** Expected Currents: 
** NormalTransistorNmos: 5.37201e+06 muA
** NormalTransistorNmos: 2.04261e+07 muA
** NormalTransistorPmos: -1.69219e+07 muA
** NormalTransistorPmos: -1.35239e+07 muA
** NormalTransistorPmos: -1.35239e+07 muA
** DiodeTransistorNmos: 1.35231e+07 muA
** DiodeTransistorNmos: 1.35231e+07 muA
** NormalTransistorNmos: 1.35231e+07 muA
** NormalTransistorNmos: 1.35231e+07 muA
** NormalTransistorPmos: -4.74779e+07 muA
** DiodeTransistorPmos: -4.74789e+07 muA
** NormalTransistorPmos: -1.35249e+07 muA
** NormalTransistorPmos: -1.35249e+07 muA
** NormalTransistorNmos: 2.2972e+08 muA
** NormalTransistorPmos: -2.29719e+08 muA
** DiodeTransistorNmos: 1.69211e+07 muA
** DiodeTransistorPmos: -5.37299e+06 muA
** NormalTransistorPmos: -5.37399e+06 muA
** DiodeTransistorPmos: -2.04269e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.06101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.634001  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outInputVoltageBiasXXpXX1: 3.40701  V
** outSourceVoltageBiasXXpXX1: 4.20301  V
** outVoltageBiasXXpXX2: 1.77601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.31901  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 2.99101  V
** sourceGCC2: 2.98601  V
** inner: 4.20301  V


.END