.suckt  two_stage_fully_differential_op_amp_60_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 outVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
m5 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m6 outFeedback outFeedback sourcePmos sourcePmos pmos
m7 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m8 FeedbackStageYinnerStageBias1 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m9 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m10 FeedbackStageYinnerStageBias2 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m11 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m15 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m16 FirstStageYsourceGCC1 outFeedback sourcePmos sourcePmos pmos
m17 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m18 FirstStageYsourceGCC2 outFeedback sourcePmos sourcePmos pmos
m19 out1FirstStage outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m20 out2FirstStage outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m21 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m22 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m23 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m24 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m25 out1 inputVoltageBiasXXnXX2 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m26 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m27 out1 outVoltageBiasXXpXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m28 SecondStage1YinnerStageBias ibias sourcePmos sourcePmos pmos
m29 out2 inputVoltageBiasXXnXX2 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m30 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m31 out2 outVoltageBiasXXpXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m32 SecondStage2YinnerStageBias ibias sourcePmos sourcePmos pmos
m33 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m34 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m35 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m36 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m37 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m38 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_60_4

