.suckt  symmetrical_op_amp129 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage out2FirstStage out1FirstStage out1FirstStage nmos
m2 out1FirstStage out1FirstStage sourceNmos sourceNmos nmos
m3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage nmos
m4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m5 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m6 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m7 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m8 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c1 out sourceNmos 
m9 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m10 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m11 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m12 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m13 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos
m14 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m15 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m17 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m18 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end symmetrical_op_amp129

