** Name: two_stage_single_output_op_amp_40_7

.MACRO two_stage_single_output_op_amp_40_7 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=49e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=34e-6
m4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=69e-6
m5 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=8e-6 W=69e-6
m6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=21e-6
m7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=36e-6
m8 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=34e-6
m9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=49e-6
m10 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=30e-6
m11 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=567e-6
m12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=36e-6
m13 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=69e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=111e-6
m15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=8e-6 W=69e-6
m16 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=37e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_40_7

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 3.45901 mW
** Area: 4823 (mu_m)^2
** Transit frequency: 2.59701 MHz
** Transit frequency with error factor: 2.595 MHz
** Slew rate: 3.98926 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** negPSRR: 97 dB
** posPSRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 0.190001 V
** VcmMax: 3.76001 V
** VcmMin: 1.37001 V


** Expected Currents: 
** NormalTransistorNmos: 2.99901e+07 muA
** NormalTransistorPmos: -5.19129e+07 muA
** DiodeTransistorPmos: -1.82099e+07 muA
** NormalTransistorPmos: -1.82089e+07 muA
** NormalTransistorPmos: -1.82099e+07 muA
** DiodeTransistorPmos: -1.82089e+07 muA
** NormalTransistorNmos: 3.64171e+07 muA
** DiodeTransistorNmos: 3.64161e+07 muA
** NormalTransistorNmos: 1.82091e+07 muA
** NormalTransistorNmos: 1.82091e+07 muA
** NormalTransistorNmos: 5.63514e+08 muA
** NormalTransistorPmos: -5.63513e+08 muA
** DiodeTransistorNmos: 5.19121e+07 muA
** NormalTransistorNmos: 5.19121e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.99909e+07 muA


** Expected Voltages: 
** ibias: 0.593001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.74701  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.12801  V
** outSourceVoltageBiasXXnXX1: 0.564001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.26501  V
** innerTransistorStack1Load1: 4.26501  V
** out1: 3.35801  V
** sourceTransconductance: 1.85001  V
** inner: 0.564001  V


.END