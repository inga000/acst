** Name: one_stage_single_output_op_amp48

.MACRO one_stage_single_output_op_amp48 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=13e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=113e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=161e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=161e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=9e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=150e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=150e-6
mFoldedCascodeFirstStageLoad9 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=9e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=161e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=354e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=354e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=95e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=107e-6
mFoldedCascodeFirstStageLoad15 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=161e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp48

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 2.06701 mW
** Area: 3868 (mu_m)^2
** Transit frequency: 5.04401 MHz
** Transit frequency with error factor: 5.04364 MHz
** Slew rate: 4.74343 V/mu_s
** Phase margin: 88.8085°
** CMRR: 138 dB
** VoutMax: 4.07001 V
** VoutMin: 1.06001 V
** VcmMax: 4.05001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.07611e+08 muA
** NormalTransistorNmos: 9.50451e+07 muA
** NormalTransistorNmos: 1.42848e+08 muA
** NormalTransistorNmos: 9.50451e+07 muA
** NormalTransistorNmos: 1.42848e+08 muA
** DiodeTransistorPmos: -9.50459e+07 muA
** NormalTransistorPmos: -9.50469e+07 muA
** NormalTransistorPmos: -9.50459e+07 muA
** DiodeTransistorPmos: -9.50469e+07 muA
** NormalTransistorPmos: -9.56069e+07 muA
** NormalTransistorPmos: -4.78029e+07 muA
** NormalTransistorPmos: -4.78029e+07 muA
** DiodeTransistorNmos: 1.07612e+08 muA
** DiodeTransistorNmos: 1.07613e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.40101  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.25401  V
** innerTransistorStack1Load2: 4.25301  V
** out1: 3.50801  V
** sourceGCC1: 0.494001  V
** sourceGCC2: 0.494001  V
** sourceTransconductance: 3.21401  V


.END