** Name: two_stage_single_output_op_amp_16_2

.MACRO two_stage_single_output_op_amp_16_2 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=21e-6
mSecondStage1StageBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=17e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=28e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=190e-6
mSimpleFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=540e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=477e-6
mSecondStage1Transconductor8 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=214e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=21e-6
mMainBias10 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=81e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=116e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=540e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=190e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=237e-6
mSecondStage1StageBias15 out ibias sourcePmos sourcePmos pmos4 L=4e-6 W=502e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=116e-6
mMainBias17 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=18e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.5e-12
.EOM two_stage_single_output_op_amp_16_2

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 2.04801 mW
** Area: 14972 (mu_m)^2
** Transit frequency: 3.92001 MHz
** Transit frequency with error factor: 3.9079 MHz
** Slew rate: 6.37856 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** negPSRR: 93 dB
** posPSRR: 110 dB
** VoutMax: 4.72001 V
** VoutMin: 0.320001 V
** VcmMax: 3.09001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 3.03011e+07 muA
** NormalTransistorPmos: -6.47199e+06 muA
** NormalTransistorPmos: -8.50509e+07 muA
** DiodeTransistorNmos: 4.25771e+07 muA
** NormalTransistorNmos: 4.25771e+07 muA
** NormalTransistorPmos: -8.51569e+07 muA
** DiodeTransistorPmos: -8.51579e+07 muA
** NormalTransistorPmos: -4.25779e+07 muA
** NormalTransistorPmos: -4.25779e+07 muA
** NormalTransistorNmos: 1.82713e+08 muA
** NormalTransistorNmos: 1.82712e+08 muA
** NormalTransistorPmos: -1.82712e+08 muA
** DiodeTransistorNmos: 6.47101e+06 muA
** DiodeTransistorNmos: 8.50501e+07 muA
** DiodeTransistorPmos: -3.03019e+07 muA
** NormalTransistorPmos: -3.03029e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.15201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.729001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.49601  V
** outSourceVoltageBiasXXpXX1: 4.24801  V
** outVoltageBiasXXnXX0: 0.616001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.559001  V
** sourceTransconductance: 3.46801  V
** innerTransconductance: 0.150001  V
** inner: 4.24801  V


.END