** Name: symmetrical_op_amp149

.MACRO symmetrical_op_amp149 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=13e-6
mMainBias3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=57e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=174e-6
mSymmetricalFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=171e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=15e-6
mSymmetricalFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=15e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=42e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=42e-6
mSymmetricalFirstStageLoad11 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=21e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor12 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=3e-6 W=52e-6
mSecondStage1Transconductor13 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=52e-6
mSymmetricalFirstStageLoad14 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=21e-6
mMainBias15 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=540e-6
mSymmetricalFirstStageStageBias16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=171e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=174e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=57e-6
mSymmetricalFirstStageTransconductor19 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=234e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=105e-6
mSymmetricalFirstStageTransconductor21 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=234e-6
mMainBias22 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=264e-6
mMainBias23 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=56e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp149

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 2.99001 mW
** Area: 13684 (mu_m)^2
** Transit frequency: 3.96701 MHz
** Transit frequency with error factor: 3.96712 MHz
** Slew rate: 4.22144 V/mu_s
** Phase margin: 83.6519°
** CMRR: 153 dB
** negPSRR: 53 dB
** posPSRR: 76 dB
** VoutMax: 4.54001 V
** VoutMin: 0.320001 V
** VcmMax: 3.26001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.06136e+08 muA
** NormalTransistorPmos: -9.89799e+06 muA
** NormalTransistorPmos: -4.69249e+07 muA
** NormalTransistorNmos: 1.52121e+07 muA
** NormalTransistorNmos: 1.52111e+07 muA
** NormalTransistorNmos: 1.52121e+07 muA
** NormalTransistorNmos: 1.52111e+07 muA
** NormalTransistorPmos: -3.04249e+07 muA
** DiodeTransistorPmos: -3.04239e+07 muA
** NormalTransistorPmos: -1.52129e+07 muA
** NormalTransistorPmos: -1.52129e+07 muA
** NormalTransistorNmos: 4.22851e+07 muA
** NormalTransistorNmos: 4.22861e+07 muA
** NormalTransistorPmos: -4.22859e+07 muA
** NormalTransistorPmos: -4.22869e+07 muA
** DiodeTransistorPmos: -4.22859e+07 muA
** NormalTransistorNmos: 4.22851e+07 muA
** NormalTransistorNmos: 4.22861e+07 muA
** DiodeTransistorNmos: 9.89701e+06 muA
** DiodeTransistorNmos: 4.69241e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -4.06135e+08 muA


** Expected Voltages: 
** ibias: 3.42601  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.560001  V
** innerComplementarySecondStage: 4.12601  V
** out: 2.5  V
** out1FirstStage: 0.560001  V
** out2FirstStage: 0.729001  V
** outSourceVoltageBiasXXpXX1: 4.21401  V
** outVoltageBiasXXnXX0: 0.616001  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.163001  V
** innerTransistorStack2Load1: 0.163001  V
** sourceTransconductance: 3.23401  V
** innerStageBias: 4.40001  V
** innerTransconductance: 0.155001  V
** inner: 0.155001  V
** inner: 4.21101  V


.END