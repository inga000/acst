.suckt  complementary_op_amp24 ibias in1 in2 out sourceNmos sourcePmos
m_Complementary_MainBias_1 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_MainBias_2 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_MainBias_3 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_4 FirstStageYinnerSourceLoadPmos outInputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m_Complementary_FirstStage_Load_5 FirstStageYinnerTransistorStack1LoadNmos outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_6 out outInputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m_Complementary_FirstStage_Load_7 FirstStageYinnerTransistorStack2LoadNmos outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_8 FirstStageYinnerSourceLoadPmos outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m_Complementary_FirstStage_Load_9 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_10 out outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m_Complementary_FirstStage_Load_11 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_StageBias_12 FirstStageYsourceTransconductanceNmos outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_Complementary_FirstStage_StageBias_13 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_14 FirstStageYsourceTransconductancePmos ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_Complementary_FirstStage_StageBias_15 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Transconductor_16 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_17 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_18 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m_Complementary_FirstStage_Transconductor_19 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c_Complementary_Load_Capacitor_1 out sourceNmos 
m_Complementary_MainBias_20 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_Complementary_MainBias_21 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_MainBias_22 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m_Complementary_MainBias_23 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_MainBias_24 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_Complementary_MainBias_25 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_MainBias_26 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end complementary_op_amp24

