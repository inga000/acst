.suckt  two_stage_fully_differential_op_amp_23_1 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 outVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m5 outFeedback outFeedback sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m7 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m8 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m9 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m10 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m12 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m13 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m14 out1FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m15 FirstStageYinnerTransistorStack1Load2 outFeedback sourcePmos sourcePmos pmos
m16 out2FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m17 FirstStageYinnerTransistorStack2Load2 outFeedback sourcePmos sourcePmos pmos
m18 sourceTransconductance ibias sourceNmos sourceNmos nmos
m19 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m20 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m21 out1 out1FirstStage sourceNmos sourceNmos nmos
m22 out1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m23 out2 out2FirstStage sourceNmos sourceNmos nmos
m24 out2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m25 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
m26 ibias ibias sourceNmos sourceNmos nmos
m27 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m28 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_23_1

