** Name: one_stage_single_output_op_amp105

.MACRO one_stage_single_output_op_amp105 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=35e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=29e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=23e-6
mMainBias5 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=12e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=35e-6
mTelescopicFirstStageLoad8 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=29e-6
mMainBias9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=20e-6
mTelescopicFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=231e-6
mTelescopicFirstStageLoad11 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=82e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=9e-6 W=185e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=9e-6 W=185e-6
mTelescopicFirstStageLoad14 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=82e-6
mMainBias15 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=582e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp105

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 1.36101 mW
** Area: 5078 (mu_m)^2
** Transit frequency: 2.84501 MHz
** Transit frequency with error factor: 2.84523 MHz
** Slew rate: 11.6889 V/mu_s
** Phase margin: 85.9437°
** CMRR: 133 dB
** VoutMax: 3.08001 V
** VoutMin: 0.760001 V
** VcmMax: 3 V
** VcmMin: 1.09001 V


** Expected Currents: 
** NormalTransistorNmos: 5.95871e+07 muA
** NormalTransistorPmos: -1.81499e+07 muA
** NormalTransistorPmos: -8.72779e+07 muA
** NormalTransistorPmos: -8.72779e+07 muA
** DiodeTransistorNmos: 8.72771e+07 muA
** DiodeTransistorNmos: 8.72761e+07 muA
** NormalTransistorNmos: 8.72771e+07 muA
** NormalTransistorNmos: 8.72761e+07 muA
** NormalTransistorPmos: -2.34142e+08 muA
** NormalTransistorPmos: -2.34143e+08 muA
** NormalTransistorPmos: -8.72769e+07 muA
** NormalTransistorPmos: -8.72769e+07 muA
** DiodeTransistorNmos: 1.81491e+07 muA
** DiodeTransistorPmos: -5.95879e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.671001  V
** outVoltageBiasXXpXX1: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.54901  V
** innerStageBias: 4.19301  V
** innerTransistorStack1Load2: 0.576001  V
** innerTransistorStack2Load2: 0.575001  V
** out1: 1.16901  V
** sourceGCC1: 2.98801  V
** sourceGCC2: 2.98801  V


.END