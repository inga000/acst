** Name: two_stage_single_output_op_amp_3_1

.MACRO two_stage_single_output_op_amp_3_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=101e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=101e-6
mSecondStage1Transconductor5 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=400e-6
mSimpleFirstStageLoad6 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=31e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=19e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=221e-6
mMainBias9 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=97e-6
mSecondStage1StageBias10 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=349e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=19e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_3_1

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 1.55601 mW
** Area: 3818 (mu_m)^2
** Transit frequency: 4.51001 MHz
** Transit frequency with error factor: 4.49323 MHz
** Slew rate: 6.19765 V/mu_s
** Phase margin: 62.4525°
** CMRR: 92 dB
** negPSRR: 94 dB
** posPSRR: 210 dB
** VoutMax: 4.84001 V
** VoutMin: 0.150001 V
** VcmMax: 3.53001 V
** VcmMin: 0.260001 V


** Expected Currents: 
** NormalTransistorPmos: -4.1875e+07 muA
** DiodeTransistorNmos: 4.82291e+07 muA
** NormalTransistorNmos: 4.82281e+07 muA
** NormalTransistorNmos: 4.82291e+07 muA
** NormalTransistorPmos: -9.64569e+07 muA
** NormalTransistorPmos: -4.82279e+07 muA
** NormalTransistorPmos: -4.82279e+07 muA
** NormalTransistorNmos: 1.52801e+08 muA
** NormalTransistorPmos: -1.528e+08 muA
** DiodeTransistorNmos: 4.18741e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.827001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.81401  V


.END