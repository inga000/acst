** Name: symmetrical_op_amp27

.MACRO symmetrical_op_amp27 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=47e-6
mSecondStage1StageBias2 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=61e-6
mSecondStage1StageBias3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
mSymmetricalFirstStageLoad4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=83e-6
mSymmetricalFirstStageLoad5 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=83e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=9e-6 W=600e-6
mMainBias7 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos4 L=9e-6 W=47e-6
mSymmetricalFirstStageTransconductor8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=44e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias9 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=61e-6
mSecondStage1StageBias10 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos4 L=1e-6 W=32e-6
mSymmetricalFirstStageTransconductor11 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=44e-6
mSecondStage1Transconductor12 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=121e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor13 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=121e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=6e-6 W=134e-6
mSecondStage1Transconductor15 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=6e-6 W=134e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp27

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 1.68601 mW
** Area: 8750 (mu_m)^2
** Transit frequency: 8.00401 MHz
** Transit frequency with error factor: 8.00436 MHz
** Slew rate: 9.43293 V/mu_s
** Phase margin: 61.3065°
** CMRR: 144 dB
** negPSRR: 51 dB
** posPSRR: 44 dB
** VoutMax: 4.31001 V
** VoutMin: 0.780001 V
** VcmMax: 4.63001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00461e+07 muA
** DiodeTransistorPmos: -6.41299e+07 muA
** DiodeTransistorPmos: -6.41299e+07 muA
** NormalTransistorNmos: 1.28258e+08 muA
** NormalTransistorNmos: 6.41291e+07 muA
** NormalTransistorNmos: 6.41291e+07 muA
** NormalTransistorNmos: 9.44931e+07 muA
** DiodeTransistorNmos: 9.44921e+07 muA
** NormalTransistorPmos: -9.44939e+07 muA
** NormalTransistorPmos: -9.44929e+07 muA
** NormalTransistorNmos: 9.44931e+07 muA
** NormalTransistorPmos: -9.44939e+07 muA
** NormalTransistorPmos: -9.44929e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.00469e+07 muA


** Expected Voltages: 
** ibias: 0.555001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 4.22801  V
** inStageBiasComplementarySecondStage: 0.596001  V
** innerComplementarySecondStage: 1.18701  V
** out: 2.5  V
** outFirstStage: 4.22801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.90901  V
** innerTransconductance: 4.73501  V
** inner: 4.73501  V


.END