.suckt  two_stage_fully_differential_op_amp_45_6 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outInputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_3 outVoltageBiasXXpXX3 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_4 outVoltageBiasXXpXX4 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_5 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_6 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_7 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_Load_8 outFeedback outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_10 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackStage_Transconductor_11 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FeedbackStage_Transconductor_14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FirstStage_Load_15 out1FirstStage outVoltageBiasXXpXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m_FullyDifferential_FirstStage_Load_16 out2FirstStage outVoltageBiasXXpXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m_FullyDifferential_FirstStage_Load_17 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m_FullyDifferential_FirstStage_Load_18 FirstStageYinnerTransistorStack1Load2 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_19 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m_FullyDifferential_FirstStage_Load_20 FirstStageYinnerTransistorStack2Load2 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_StageBias_21 sourceTransconductance outVoltageBiasXXpXX4 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m_FullyDifferential_FirstStage_StageBias_22 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Transconductor_23 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m_FullyDifferential_FirstStage_Transconductor_24 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_Transconductor_25 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m_FullyDifferential_SecondStage1_Transconductor_26 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_27 out1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_FullyDifferential_SecondStage1_StageBias_28 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_Transconductor_29 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m_FullyDifferential_SecondStage2_Transconductor_30 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_StageBias_31 out2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m_FullyDifferential_SecondStage2_StageBias_32 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_33 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_34 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_35 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_FullyDifferential_MainBias_36 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_37 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m_FullyDifferential_MainBias_38 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_39 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourceTransconductance sourceTransconductance pmos
m_FullyDifferential_MainBias_40 outVoltageBiasXXpXX4 outVoltageBiasXXpXX4 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_41 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_45_6

