** Name: two_stage_single_output_op_amp_52_1

.MACRO two_stage_single_output_op_amp_52_1 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=160e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=16e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=22e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=160e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=241e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=241e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=6e-6 W=237e-6
mMainBias10 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=43e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=425e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=219e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=144e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=409e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=185e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=185e-6
mMainBias17 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=75e-6
mSecondStage1StageBias18 out inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=592e-6
mFoldedCascodeFirstStageLoad19 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=409e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.6001e-12
.EOM two_stage_single_output_op_amp_52_1

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 7.75601 mW
** Area: 10471 (mu_m)^2
** Transit frequency: 12.2881 MHz
** Transit frequency with error factor: 12.2877 MHz
** Slew rate: 12.0666 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 4.61001 V
** VoutMin: 0.150001 V
** VcmMax: 5.02001 V
** VcmMin: 0.790001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorNmos: 3.01991e+07 muA
** NormalTransistorPmos: -1.01588e+08 muA
** NormalTransistorPmos: -1.66108e+08 muA
** NormalTransistorPmos: -2.49165e+08 muA
** NormalTransistorPmos: -1.66108e+08 muA
** NormalTransistorPmos: -2.49165e+08 muA
** DiodeTransistorNmos: 1.66109e+08 muA
** NormalTransistorNmos: 1.66109e+08 muA
** NormalTransistorNmos: 1.66109e+08 muA
** NormalTransistorNmos: 1.66113e+08 muA
** NormalTransistorNmos: 8.30561e+07 muA
** NormalTransistorNmos: 8.30561e+07 muA
** NormalTransistorNmos: 8.09467e+08 muA
** NormalTransistorPmos: -8.09466e+08 muA
** DiodeTransistorNmos: 1.01589e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -3.01999e+07 muA


** Expected Voltages: 
** ibias: 0.629001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.950001  V
** inputVoltageBiasXXpXX2: 4.04601  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.356001  V
** out1: 0.561001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.93801  V


.END