** Name: two_stage_single_output_op_amp_29_7

.MACRO two_stage_single_output_op_amp_29_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=13e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=250e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=13e-6
mSimpleFirstStageStageBias5 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=387e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=31e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=464e-6
mSecondStage1StageBias8 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=469e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=31e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=16e-6
mMainBias11 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=31e-6
mSecondStage1Transconductor12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=250e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_29_7

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 3.55501 mW
** Area: 8001 (mu_m)^2
** Transit frequency: 6.84201 MHz
** Transit frequency with error factor: 6.79842 MHz
** Slew rate: 12.371 V/mu_s
** Phase margin: 60.1606°
** CMRR: 87 dB
** negPSRR: 127 dB
** posPSRR: 85 dB
** VoutMax: 4.82001 V
** VoutMin: 0.210001 V
** VcmMax: 4.66001 V
** VcmMin: 1.92001 V


** Expected Currents: 
** NormalTransistorNmos: 1.24131e+07 muA
** NormalTransistorPmos: -2.94519e+07 muA
** DiodeTransistorPmos: -1.48193e+08 muA
** NormalTransistorPmos: -1.48193e+08 muA
** NormalTransistorNmos: 2.96386e+08 muA
** NormalTransistorNmos: 2.96385e+08 muA
** NormalTransistorNmos: 1.48194e+08 muA
** NormalTransistorNmos: 1.48194e+08 muA
** NormalTransistorNmos: 3.62695e+08 muA
** NormalTransistorPmos: -3.62694e+08 muA
** DiodeTransistorNmos: 2.94511e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.24139e+07 muA


** Expected Voltages: 
** ibias: 0.618001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.768001  V
** out: 2.5  V
** outFirstStage: 4.25301  V
** outVoltageBiasXXpXX0: 3.70401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.213001  V
** out1: 4.25301  V
** sourceTransconductance: 1.34501  V


.END