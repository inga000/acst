** Name: two_stage_single_output_op_amp_10_11

.MACRO two_stage_single_output_op_amp_10_11 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=21e-6
m3 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=213e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=48e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=514e-6
m6 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=38e-6
m7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
m8 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=217e-6
m9 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=341e-6
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
m11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=86e-6
m12 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=549e-6
m13 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=514e-6
m14 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=40e-6
m15 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=561e-6
m16 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=514e-6
m17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=206e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.20001e-12
.EOM two_stage_single_output_op_amp_10_11

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 12.5341 mW
** Area: 9733 (mu_m)^2
** Transit frequency: 7.32301 MHz
** Transit frequency with error factor: 7.30972 MHz
** Slew rate: 19.4246 V/mu_s
** Phase margin: 60.1606°
** CMRR: 100 dB
** negPSRR: 145 dB
** posPSRR: 93 dB
** VoutMax: 4.25 V
** VoutMin: 0.670001 V
** VcmMax: 4.39001 V
** VcmMin: 1.01001 V


** Expected Currents: 
** NormalTransistorNmos: 3.08965e+08 muA
** NormalTransistorNmos: 4.87363e+08 muA
** NormalTransistorPmos: -7.99549e+08 muA
** DiodeTransistorPmos: -6.03469e+07 muA
** NormalTransistorPmos: -6.03469e+07 muA
** NormalTransistorPmos: -6.03469e+07 muA
** NormalTransistorNmos: 1.20693e+08 muA
** NormalTransistorNmos: 6.03461e+07 muA
** NormalTransistorNmos: 6.03461e+07 muA
** NormalTransistorNmos: 7.80276e+08 muA
** NormalTransistorNmos: 7.80275e+08 muA
** NormalTransistorPmos: -7.80275e+08 muA
** NormalTransistorPmos: -7.80276e+08 muA
** DiodeTransistorNmos: 7.9955e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.08964e+08 muA
** DiodeTransistorPmos: -4.87362e+08 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.97601  V
** outVoltageBiasXXnXX1: 1.07901  V
** outVoltageBiasXXpXX0: 3.94501  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.54001  V
** out1: 4.27401  V
** sourceTransconductance: 1.67101  V
** innerStageBias: 0.183001  V
** innerTransconductance: 4.54001  V


.END