.suckt  two_stage_single_output_op_amp_39_7 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mMainBias2 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad5 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos
mSecondStage1Transconductor12 out outFirstStage sourcePmos sourcePmos pmos
mMainBias13 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias14 ibias ibias sourceNmos sourceNmos nmos
mMainBias15 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_39_7

