** Name: two_stage_single_output_op_amp_35_9

.MACRO two_stage_single_output_op_amp_35_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=29e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=8e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=134e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=141e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=7e-6 W=63e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=14e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=51e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=31e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=29e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=36e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=134e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=31e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=141e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=473e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=7e-6 W=63e-6
mMainBias18 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=43e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_35_9

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 3.36701 mW
** Area: 10702 (mu_m)^2
** Transit frequency: 3.25301 MHz
** Transit frequency with error factor: 3.2508 MHz
** Slew rate: 3.60224 V/mu_s
** Phase margin: 64.7443°
** CMRR: 105 dB
** negPSRR: 97 dB
** posPSRR: 93 dB
** VoutMax: 4.25 V
** VoutMin: 1.70001 V
** VcmMax: 3.90001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 1.16761e+07 muA
** NormalTransistorPmos: -3.51939e+07 muA
** DiodeTransistorPmos: -8.15099e+06 muA
** DiodeTransistorPmos: -8.15199e+06 muA
** NormalTransistorPmos: -8.15299e+06 muA
** NormalTransistorPmos: -8.15199e+06 muA
** NormalTransistorNmos: 1.63031e+07 muA
** NormalTransistorNmos: 1.63021e+07 muA
** NormalTransistorNmos: 8.15201e+06 muA
** NormalTransistorNmos: 8.15201e+06 muA
** NormalTransistorNmos: 6.0032e+08 muA
** DiodeTransistorNmos: 6.00319e+08 muA
** NormalTransistorPmos: -6.00319e+08 muA
** DiodeTransistorNmos: 3.51931e+07 muA
** NormalTransistorNmos: 3.51931e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.16769e+07 muA


** Expected Voltages: 
** ibias: 1.11701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.13201  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 2.10601  V
** outSourceVoltageBiasXXnXX1: 1.05301  V
** outSourceVoltageBiasXXnXX2: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.28601  V
** innerStageBias: 0.512001  V
** innerTransistorStack2Load1: 4.28701  V
** out1: 3.49801  V
** sourceTransconductance: 1.91801  V
** inner: 1.05301  V


.END