.suckt  one_stage_single_output_op_amp164 ibias in1 in2 out sourceNmos sourcePmos
m_SingleOutput_MainBias_1 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_4 out outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_6 FirstStageYout1 ibias sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_7 out ibias sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_StageBias_8 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_SingleOutput_FirstStage_StageBias_9 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Transconductor_10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_SingleOutput_FirstStage_Transconductor_11 out in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_SingleOutput_Load_Capacitor_1 out sourceNmos 
m_SingleOutput_MainBias_12 ibias ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_13 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_SingleOutput_MainBias_14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_15 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end one_stage_single_output_op_amp164

