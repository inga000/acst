** Name: one_stage_single_output_op_amp79

.MACRO one_stage_single_output_op_amp79 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=21e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=118e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=117e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=117e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=261e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=72e-6
mFoldedCascodeFirstStageLoad12 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=261e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=361e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=343e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=343e-6
mFoldedCascodeFirstStageLoad16 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=361e-6
mMainBias17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
mMainBias18 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp79

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 3.91101 mW
** Area: 5275 (mu_m)^2
** Transit frequency: 9.90101 MHz
** Transit frequency with error factor: 9.90077 MHz
** Slew rate: 11.5102 V/mu_s
** Phase margin: 87.0896°
** CMRR: 138 dB
** VoutMax: 4.01001 V
** VoutMin: 0.540001 V
** VcmMax: 5.17001 V
** VcmMin: 1.54001 V


** Expected Currents: 
** NormalTransistorPmos: -4.66379e+07 muA
** NormalTransistorPmos: -2.00159e+07 muA
** NormalTransistorPmos: -2.31838e+08 muA
** NormalTransistorPmos: -3.47756e+08 muA
** NormalTransistorPmos: -2.31841e+08 muA
** NormalTransistorPmos: -3.47759e+08 muA
** NormalTransistorNmos: 2.3184e+08 muA
** NormalTransistorNmos: 2.31841e+08 muA
** NormalTransistorNmos: 2.31842e+08 muA
** NormalTransistorNmos: 2.31841e+08 muA
** NormalTransistorNmos: 2.31838e+08 muA
** NormalTransistorNmos: 2.31837e+08 muA
** NormalTransistorNmos: 1.1592e+08 muA
** NormalTransistorNmos: 1.1592e+08 muA
** DiodeTransistorNmos: 4.66371e+07 muA
** DiodeTransistorNmos: 2.00151e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.15001  V
** outVoltageBiasXXnXX2: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.353001  V
** innerTransistorStack1Load2: 0.540001  V
** innerTransistorStack2Load2: 0.541001  V
** out1: 0.746001  V
** sourceGCC1: 4.22401  V
** sourceGCC2: 4.22401  V
** sourceTransconductance: 1.91001  V


.END