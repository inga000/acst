.suckt  two_stage_fully_differential_op_amp_44_5 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 outInputVoltageBiasXXpXX3 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m4 outVoltageBiasXXpXX4 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m5 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX5 sourcePmos sourcePmos pmos
m6 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m7 outFeedback outFeedback sourceNmos sourceNmos nmos
m8 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m9 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXpXX5 sourcePmos sourcePmos pmos
m10 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m11 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXpXX5 sourcePmos sourcePmos pmos
m12 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m13 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m14 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m15 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m16 out1FirstStage outVoltageBiasXXpXX4 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m17 out2FirstStage outVoltageBiasXXpXX4 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m18 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m19 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m20 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m21 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m22 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m23 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m24 out1 out1FirstStage sourceNmos sourceNmos nmos
m25 out1 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m26 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m27 out2 out2FirstStage sourceNmos sourceNmos nmos
m28 out2 outInputVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos
m29 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m30 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m31 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m32 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m33 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m34 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m35 outInputVoltageBiasXXpXX3 outInputVoltageBiasXXpXX3 VoltageBiasXXpXX3Yinner VoltageBiasXXpXX3Yinner pmos
m36 VoltageBiasXXpXX3Yinner outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m37 outVoltageBiasXXpXX4 outVoltageBiasXXpXX4 sourceTransconductance sourceTransconductance pmos
m38 ibias ibias outSourceVoltageBiasXXpXX5 outSourceVoltageBiasXXpXX5 pmos
m39 outSourceVoltageBiasXXpXX5 outSourceVoltageBiasXXpXX5 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_44_5

