** Name: two_stage_single_output_op_amp_52_7

.MACRO two_stage_single_output_op_amp_52_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=15e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=44e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=33e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=15e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=29e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=29e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=13e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=594e-6
mFoldedCascodeFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=54e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=45e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=580e-6
mFoldedCascodeFirstStageLoad16 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=45e-6
mMainBias17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=292e-6
mMainBias18 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_52_7

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 6.28301 mW
** Area: 7135 (mu_m)^2
** Transit frequency: 3.72301 MHz
** Transit frequency with error factor: 3.72291 MHz
** Slew rate: 4.03358 V/mu_s
** Phase margin: 67.6091°
** CMRR: 141 dB
** VoutMax: 4.25 V
** VoutMin: 0.180001 V
** VcmMax: 5.17001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorPmos: -2.9432e+08 muA
** NormalTransistorPmos: -4.63129e+07 muA
** NormalTransistorPmos: -1.825e+07 muA
** NormalTransistorPmos: -2.73739e+07 muA
** NormalTransistorPmos: -1.825e+07 muA
** NormalTransistorPmos: -2.73739e+07 muA
** DiodeTransistorNmos: 1.82491e+07 muA
** NormalTransistorNmos: 1.82491e+07 muA
** NormalTransistorNmos: 1.82491e+07 muA
** NormalTransistorNmos: 1.82491e+07 muA
** NormalTransistorNmos: 9.12501e+06 muA
** NormalTransistorNmos: 9.12501e+06 muA
** NormalTransistorNmos: 8.41282e+08 muA
** NormalTransistorPmos: -8.41281e+08 muA
** DiodeTransistorNmos: 2.94321e+08 muA
** DiodeTransistorNmos: 4.63121e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.09701  V
** outVoltageBiasXXnXX2: 0.588001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.538001  V
** out1: 0.743001  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.92201  V


.END