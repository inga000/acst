.suckt  two_stage_fully_differential_op_amp_27_7 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m4 outFeedback outFeedback sourceNmos sourceNmos nmos
m5 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m7 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m8 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m9 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m10 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m11 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m12 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m13 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m14 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m15 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m16 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m17 out1 ibias sourceNmos sourceNmos nmos
m18 out1 out1FirstStage sourcePmos sourcePmos pmos
m19 out2 ibias sourceNmos sourceNmos nmos
m20 out2 out2FirstStage sourcePmos sourcePmos pmos
m21 ibias ibias sourceNmos sourceNmos nmos
m22 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m24 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_27_7

