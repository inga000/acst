** Name: two_stage_single_output_op_amp_129_4

.MACRO two_stage_single_output_op_amp_129_4 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=28e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=148e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
m5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=189e-6
m6 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=166e-6
m7 outFirstStage outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=429e-6
m8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=278e-6
m9 FirstStageYout1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=429e-6
m10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=500e-6
m11 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=600e-6
m12 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=479e-6
m13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=292e-6
m14 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=402e-6
m15 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=533e-6
m16 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=2e-6 W=189e-6
m17 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=292e-6
m18 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=220e-6
m19 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=598e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 19.7001e-12
.EOM two_stage_single_output_op_amp_129_4

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 14.9991 mW
** Area: 14749 (mu_m)^2
** Transit frequency: 3.33201 MHz
** Transit frequency with error factor: 3.29875 MHz
** Slew rate: 5.87857 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.53001 V
** VoutMin: 0.300001 V
** VcmMax: 3.86001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 5.31703e+08 muA
** NormalTransistorPmos: -2.12617e+08 muA
** NormalTransistorPmos: -2.81885e+08 muA
** NormalTransistorPmos: -7.5831e+08 muA
** NormalTransistorPmos: -7.5831e+08 muA
** DiodeTransistorPmos: -7.5831e+08 muA
** NormalTransistorNmos: 8.17086e+08 muA
** NormalTransistorNmos: 8.17086e+08 muA
** NormalTransistorPmos: -1.17549e+08 muA
** NormalTransistorPmos: -5.87749e+07 muA
** NormalTransistorPmos: -5.87749e+07 muA
** NormalTransistorNmos: 3.19521e+08 muA
** NormalTransistorNmos: 3.1952e+08 muA
** NormalTransistorPmos: -3.1952e+08 muA
** NormalTransistorPmos: -3.19521e+08 muA
** DiodeTransistorNmos: 2.12618e+08 muA
** DiodeTransistorNmos: 2.81886e+08 muA
** DiodeTransistorPmos: -5.31702e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX1: 0.706001  V
** outVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 3.76301  V
** out1: 2.77601  V
** sourceTransconductance: 3.34401  V
** innerStageBias: 4.42201  V
** innerTransconductance: 0.150001  V


.END