** Name: two_stage_single_output_op_amp_114_8

.MACRO two_stage_single_output_op_amp_114_8 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=23e-6
m2 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=2e-6 W=5e-6
m3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=137e-6
m4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=46e-6
m5 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
m6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=210e-6
m7 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=44e-6
m8 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=44e-6
m9 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=544e-6
m10 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=8e-6 W=27e-6
m11 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=46e-6
m12 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=8e-6 W=27e-6
m13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=27e-6
m14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=8e-6 W=27e-6
m15 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=527e-6
m16 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=137e-6
m17 inputVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=107e-6
m18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=533e-6
m19 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=44e-6
m20 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=497e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_114_8

** Expected Performance Values: 
** Gain: 103 dB
** Power consumption: 3.54001 mW
** Area: 9291 (mu_m)^2
** Transit frequency: 3.01901 MHz
** Transit frequency with error factor: 3.01862 MHz
** Slew rate: 7.64554 V/mu_s
** Phase margin: 69.9009°
** CMRR: 96 dB
** VoutMax: 4.77001 V
** VoutMin: 0.710001 V
** VcmMax: 4.47001 V
** VcmMin: 1.52001 V


** Expected Currents: 
** NormalTransistorNmos: 4.32131e+07 muA
** NormalTransistorPmos: -1.02274e+08 muA
** NormalTransistorPmos: -2.16879e+07 muA
** NormalTransistorNmos: 6.42901e+06 muA
** NormalTransistorNmos: 6.42901e+06 muA
** DiodeTransistorPmos: -6.42999e+06 muA
** NormalTransistorPmos: -6.42999e+06 muA
** NormalTransistorNmos: 3.45441e+07 muA
** DiodeTransistorNmos: 3.45431e+07 muA
** NormalTransistorNmos: 6.42901e+06 muA
** NormalTransistorNmos: 6.42901e+06 muA
** NormalTransistorNmos: 5.1806e+08 muA
** NormalTransistorNmos: 5.18059e+08 muA
** NormalTransistorPmos: -5.18059e+08 muA
** DiodeTransistorNmos: 1.02275e+08 muA
** NormalTransistorNmos: 1.02274e+08 muA
** DiodeTransistorNmos: 2.16871e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -4.32139e+07 muA


** Expected Voltages: 
** ibias: 1.18001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 2.65001  V
** inputVoltageBiasXXpXX0: 4.28501  V
** out: 2.5  V
** outFirstStage: 4.20201  V
** outInputVoltageBiasXXnXX1: 1.37401  V
** outSourceVoltageBiasXXnXX1: 0.687001  V
** outSourceVoltageBiasXXnXX3: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.21401  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.625  V
** inner: 0.686001  V


.END