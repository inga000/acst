** Name: two_stage_single_output_op_amp_82_8

.MACRO two_stage_single_output_op_amp_82_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=2e-6 W=97e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=97e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=5e-6
mMainBias4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=19e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=54e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=2e-6 W=97e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=32e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=32e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=54e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=596e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=370e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=97e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=257e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=157e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=157e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=519e-6
mFoldedCascodeFirstStageLoad21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=257e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias23 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=68e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.5e-12
.EOM two_stage_single_output_op_amp_82_8

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 14.9981 mW
** Area: 4223 (mu_m)^2
** Transit frequency: 11.4151 MHz
** Transit frequency with error factor: 11.4145 MHz
** Slew rate: 13.7389 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 0.920001 V
** VcmMax: 5.17001 V
** VcmMin: 1.55001 V


** Expected Currents: 
** NormalTransistorPmos: -1.01379e+07 muA
** NormalTransistorPmos: -6.84929e+07 muA
** NormalTransistorPmos: -1.04376e+08 muA
** NormalTransistorPmos: -1.59177e+08 muA
** NormalTransistorPmos: -1.04376e+08 muA
** NormalTransistorPmos: -1.59177e+08 muA
** DiodeTransistorNmos: 1.04377e+08 muA
** NormalTransistorNmos: 1.04376e+08 muA
** NormalTransistorNmos: 1.04377e+08 muA
** DiodeTransistorNmos: 1.04376e+08 muA
** NormalTransistorNmos: 1.096e+08 muA
** DiodeTransistorNmos: 1.09599e+08 muA
** NormalTransistorNmos: 5.48001e+07 muA
** NormalTransistorNmos: 5.48001e+07 muA
** NormalTransistorNmos: 2.58267e+09 muA
** NormalTransistorNmos: 2.58267e+09 muA
** NormalTransistorPmos: -2.58266e+09 muA
** DiodeTransistorNmos: 1.01371e+07 muA
** NormalTransistorNmos: 1.01361e+07 muA
** DiodeTransistorNmos: 6.84921e+07 muA
** DiodeTransistorNmos: 6.84931e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.34401  V
** outInputVoltageBiasXXnXX2: 1.24201  V
** outSourceVoltageBiasXXnXX1: 0.672001  V
** outSourceVoltageBiasXXnXX2: 0.631001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.563001  V
** innerTransistorStack2Load2: 0.564001  V
** out1: 1.12801  V
** sourceGCC1: 4.11201  V
** sourceGCC2: 4.11201  V
** sourceTransconductance: 1.89301  V
** innerStageBias: 0.549001  V
** inner: 0.670001  V


.END