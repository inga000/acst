** Name: two_stage_single_output_op_amp_45_2

.MACRO two_stage_single_output_op_amp_45_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=55e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=487e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=50e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=101e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=157e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=157e-6
mSecondStage1Transconductor9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=328e-6
mMainBias10 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=44e-6
mSecondStage1Transconductor11 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=132e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=101e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=487e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=30e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=30e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=499e-6
mMainBias17 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=597e-6
mSecondStage1StageBias18 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=599e-6
mFoldedCascodeFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=600e-6
mMainBias20 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=252e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.7001e-12
.EOM two_stage_single_output_op_amp_45_2

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 6.56001 mW
** Area: 9682 (mu_m)^2
** Transit frequency: 4.51901 MHz
** Transit frequency with error factor: 4.51851 MHz
** Slew rate: 7.94764 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** VoutMax: 4.85001 V
** VoutMin: 0.320001 V
** VcmMax: 3.66001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 8.38041e+07 muA
** NormalTransistorPmos: -2.52257e+08 muA
** NormalTransistorPmos: -1.04755e+08 muA
** NormalTransistorNmos: 1.93602e+08 muA
** NormalTransistorNmos: 2.99028e+08 muA
** NormalTransistorNmos: 1.93602e+08 muA
** NormalTransistorNmos: 2.99028e+08 muA
** DiodeTransistorPmos: -1.93601e+08 muA
** NormalTransistorPmos: -1.93601e+08 muA
** NormalTransistorPmos: -1.93601e+08 muA
** NormalTransistorPmos: -2.10848e+08 muA
** NormalTransistorPmos: -1.05424e+08 muA
** NormalTransistorPmos: -1.05424e+08 muA
** NormalTransistorNmos: 2.53103e+08 muA
** NormalTransistorNmos: 2.53102e+08 muA
** NormalTransistorPmos: -2.53102e+08 muA
** DiodeTransistorNmos: 2.52258e+08 muA
** DiodeTransistorNmos: 1.04756e+08 muA
** DiodeTransistorPmos: -8.38049e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.905001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.570001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.57801  V
** out1: 4.22501  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.68801  V
** innerTransconductance: 0.349001  V


.END