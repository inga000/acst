.suckt  two_stage_single_output_op_amp_121_2 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 outVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
m5 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m6 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m7 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m8 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos
m9 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m10 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos
m11 sourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m12 FirstStageYinnerStageBias outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c2 out sourceNmos 
m15 out inputVoltageBiasXXnXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m16 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m17 out ibias sourcePmos sourcePmos pmos
m18 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
m19 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m20 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m21 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m22 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_121_2

