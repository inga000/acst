** Name: two_stage_single_output_op_amp_107_7

.MACRO two_stage_single_output_op_amp_107_7 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=32e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=10e-6
m4 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
m5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=193e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=470e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=37e-6
m8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
m9 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=37e-6
m10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=43e-6
m11 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=43e-6
m12 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=20e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=188e-6
m14 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=5e-6 W=74e-6
m15 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=28e-6
m16 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=599e-6
m17 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=5e-6 W=74e-6
m18 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=82e-6
m19 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=119e-6
m20 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=119e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.80001e-12
.EOM two_stage_single_output_op_amp_107_7

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 14.9961 mW
** Area: 7542 (mu_m)^2
** Transit frequency: 2.78401 MHz
** Transit frequency with error factor: 2.78431 MHz
** Slew rate: 24.449 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 3 V
** VoutMin: 0.260001 V
** VcmMax: 3.03001 V
** VcmMin: -0.199999 V


** Expected Currents: 
** NormalTransistorNmos: 1.43482e+08 muA
** NormalTransistorPmos: -4.07259e+07 muA
** NormalTransistorPmos: -5.66579e+07 muA
** NormalTransistorPmos: -1.17469e+07 muA
** NormalTransistorPmos: -1.17469e+07 muA
** NormalTransistorNmos: 1.17461e+07 muA
** NormalTransistorNmos: 1.17451e+07 muA
** NormalTransistorNmos: 1.17461e+07 muA
** NormalTransistorNmos: 1.17451e+07 muA
** NormalTransistorPmos: -1.66978e+08 muA
** NormalTransistorPmos: -1.66977e+08 muA
** NormalTransistorPmos: -1.17479e+07 muA
** NormalTransistorPmos: -1.17479e+07 muA
** NormalTransistorNmos: 2.7148e+09 muA
** NormalTransistorPmos: -2.71479e+09 muA
** DiodeTransistorNmos: 4.07251e+07 muA
** DiodeTransistorNmos: 5.66571e+07 muA
** DiodeTransistorPmos: -1.43481e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.06101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 2.43601  V
** outSourceVoltageBiasXXpXX2: 3.96101  V
** outVoltageBiasXXnXX2: 0.665001  V
** outVoltageBiasXXpXX1: 2.24101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.26001  V
** innerSourceLoad2: 0.555001  V
** innerStageBias: 3.80101  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 3.01601  V
** sourceGCC2: 3.01501  V


.END