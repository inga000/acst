** Name: two_stage_single_output_op_amp_1_1

.MACRO two_stage_single_output_op_amp_1_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=44e-6
mMainBias2 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSecondStage1Transconductor3 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=94e-6
mSimpleFirstStageLoad4 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=44e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=25e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=61e-6
mSecondStage1StageBias7 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=99e-6
mSimpleFirstStageTransconductor8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=25e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_1_1

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 0.832001 mW
** Area: 1073 (mu_m)^2
** Transit frequency: 2.63101 MHz
** Transit frequency with error factor: 2.61303 MHz
** Slew rate: 3.67206 V/mu_s
** Phase margin: 63.0254°
** CMRR: 87 dB
** negPSRR: 89 dB
** posPSRR: 207 dB
** VoutMax: 4.77001 V
** VoutMin: 0.150001 V
** VcmMax: 3.46001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** DiodeTransistorNmos: 2.81181e+07 muA
** NormalTransistorNmos: 2.81181e+07 muA
** NormalTransistorPmos: -5.62379e+07 muA
** NormalTransistorPmos: -2.81189e+07 muA
** NormalTransistorPmos: -2.81189e+07 muA
** NormalTransistorNmos: 9.01101e+07 muA
** NormalTransistorPmos: -9.01109e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceTransconductance: 3.81301  V


.END