.suckt  two_stage_single_output_op_amp_144_3 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad3 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad5 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad7 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias13 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mSecondStage1StageBias14 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mMainBias15 ibias ibias sourceNmos sourceNmos nmos
mMainBias16 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mMainBias17 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_144_3

