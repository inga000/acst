** Name: two_stage_single_output_op_amp_44_3

.MACRO two_stage_single_output_op_amp_44_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=11e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=127e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=106e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=14e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=66e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=66e-6
mMainBias9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=291e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=161e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=14e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=316e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=127e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=34e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=34e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=577e-6
mSecondStage1StageBias18 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=471e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=29e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_44_3

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 4.71601 mW
** Area: 7508 (mu_m)^2
** Transit frequency: 3.56801 MHz
** Transit frequency with error factor: 3.56771 MHz
** Slew rate: 3.70917 V/mu_s
** Phase margin: 66.4632°
** CMRR: 142 dB
** VoutMax: 4.47001 V
** VoutMin: 0.580001 V
** VcmMax: 4.02001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.11687e+08 muA
** NormalTransistorNmos: 1.20543e+08 muA
** NormalTransistorNmos: 1.67301e+07 muA
** NormalTransistorNmos: 2.51421e+07 muA
** NormalTransistorNmos: 1.67301e+07 muA
** NormalTransistorNmos: 2.51421e+07 muA
** NormalTransistorPmos: -1.67309e+07 muA
** NormalTransistorPmos: -1.67309e+07 muA
** DiodeTransistorPmos: -1.67309e+07 muA
** NormalTransistorPmos: -1.68269e+07 muA
** NormalTransistorPmos: -8.41299e+06 muA
** NormalTransistorPmos: -8.41299e+06 muA
** NormalTransistorNmos: 6.50709e+08 muA
** NormalTransistorPmos: -6.50708e+08 muA
** NormalTransistorPmos: -6.50709e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.11686e+08 muA
** DiodeTransistorPmos: -1.20542e+08 muA


** Expected Voltages: 
** ibias: 1.19101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.986001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX2: 4.18501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.26401  V
** out1: 3.52001  V
** sourceGCC1: 0.519001  V
** sourceGCC2: 0.519001  V
** sourceTransconductance: 3.23001  V
** innerStageBias: 4.52701  V


.END