** Name: symmetrical_op_amp8

.MACRO symmetrical_op_amp8 ibias in1 in2 out sourceNmos sourcePmos
m1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
m2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=48e-6
m3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=48e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=35e-6
m5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
m6 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=10e-6
m7 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=3e-6 W=56e-6
m8 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=56e-6
m9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=59e-6
m10 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=59e-6
m11 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=4e-6 W=44e-6
m12 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=129e-6
m13 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=135e-6
m14 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=129e-6
m15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=317e-6
m16 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp8

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 1.18701 mW
** Area: 3095 (mu_m)^2
** Transit frequency: 4.50101 MHz
** Transit frequency with error factor: 4.50148 MHz
** Slew rate: 5.60603 V/mu_s
** Phase margin: 85.3708°
** CMRR: 152 dB
** negPSRR: 50 dB
** posPSRR: 63 dB
** VoutMax: 3.99001 V
** VoutMin: 0.340001 V
** VcmMax: 3.98001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorPmos: -1.28099e+07 muA
** DiodeTransistorNmos: 4.61441e+07 muA
** DiodeTransistorNmos: 4.61441e+07 muA
** NormalTransistorPmos: -9.22899e+07 muA
** NormalTransistorPmos: -4.61449e+07 muA
** NormalTransistorPmos: -4.61449e+07 muA
** NormalTransistorNmos: 5.61861e+07 muA
** NormalTransistorNmos: 5.61871e+07 muA
** NormalTransistorPmos: -5.61869e+07 muA
** NormalTransistorPmos: -5.61879e+07 muA
** DiodeTransistorPmos: -5.61889e+07 muA
** DiodeTransistorPmos: -5.61899e+07 muA
** NormalTransistorNmos: 5.61881e+07 muA
** NormalTransistorNmos: 5.61871e+07 muA
** DiodeTransistorNmos: 1.28091e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18201  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.743001  V
** inSourceStageBiasComplementarySecondStage: 4.14401  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 3.01701  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.26401  V
** innerStageBias: 3.73301  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END