.suckt  symmetrical_op_amp98 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage ibias sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad2 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mSymmetricalFirstStageLoad3 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageLoad4 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mSymmetricalFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSymmetricalFirstStageTransconductor7 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSymmetricalFirstStageTransconductor8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1Transconductor9 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mSecondStage1Transconductor10 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias11 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos
mSecondStage1StageBias12 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias13 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias14 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mMainBias17 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos
mMainBias18 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp98

