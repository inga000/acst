.suckt  two_stage_fully_differential_op_amp_65_9 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m3 outInputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m4 outVoltageBiasXXnXX3 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m5 outVoltageBiasXXnXX4 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m6 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m7 outFeedback outFeedback sourcePmos sourcePmos pmos
m8 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m9 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m14 out1FirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m15 out2FirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m16 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m17 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m18 sourceTransconductance outVoltageBiasXXnXX4 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m19 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m20 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m21 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m22 out1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m23 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m24 out1 out1FirstStage sourcePmos sourcePmos pmos
m25 out2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m26 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m27 out2 out2FirstStage sourcePmos sourcePmos pmos
m28 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m29 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m30 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
m31 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m32 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos
m33 outVoltageBiasXXnXX4 outVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m34 ibias ibias sourceNmos sourceNmos nmos
m35 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_65_9

