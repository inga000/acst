** Name: two_stage_single_output_op_amp_19_3

.MACRO two_stage_single_output_op_amp_19_3 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=146e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=15e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=146e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=330e-6
mSimpleFirstStageLoad7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=46e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=17e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=79e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=60e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=317e-6
mMainBias12 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=68e-6
mSecondStage1StageBias13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=273e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=17e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_19_3

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 2.42901 mW
** Area: 4022 (mu_m)^2
** Transit frequency: 7.76501 MHz
** Transit frequency with error factor: 7.75365 MHz
** Slew rate: 12.8627 V/mu_s
** Phase margin: 67.0361°
** CMRR: 99 dB
** negPSRR: 100 dB
** posPSRR: 215 dB
** VoutMax: 3.95001 V
** VoutMin: 0.150001 V
** VcmMax: 3 V
** VcmMin: 0.240001 V


** Expected Currents: 
** NormalTransistorPmos: -6.89429e+07 muA
** DiodeTransistorNmos: 4.00481e+07 muA
** NormalTransistorNmos: 4.00481e+07 muA
** NormalTransistorNmos: 4.00481e+07 muA
** NormalTransistorPmos: -8.00969e+07 muA
** NormalTransistorPmos: -8.00959e+07 muA
** NormalTransistorPmos: -4.00489e+07 muA
** NormalTransistorPmos: -4.00489e+07 muA
** NormalTransistorNmos: 3.16826e+08 muA
** NormalTransistorPmos: -3.16825e+08 muA
** NormalTransistorPmos: -3.16826e+08 muA
** DiodeTransistorNmos: 6.89421e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.44101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.803001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerStageBias: 4.27701  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.42601  V
** innerStageBias: 4.25901  V


.END