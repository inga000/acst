** Name: two_stage_single_output_op_amp_5_1

.MACRO two_stage_single_output_op_amp_5_1 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m2 ibias ibias sourcePmos sourcePmos pmos4 L=8e-6 W=38e-6
m3 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=95e-6
m4 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=31e-6
m5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=31e-6
m6 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=31e-6
m7 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=31e-6
m8 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=71e-6
m9 out ibias sourcePmos sourcePmos pmos4 L=8e-6 W=346e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=21e-6
m11 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=21e-6
m12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=8e-6 W=222e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_5_1

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 0.945001 mW
** Area: 6158 (mu_m)^2
** Transit frequency: 2.81001 MHz
** Transit frequency with error factor: 2.7987 MHz
** Slew rate: 3.69374 V/mu_s
** Phase margin: 61.3065°
** CMRR: 93 dB
** negPSRR: 94 dB
** posPSRR: 198 dB
** VoutMax: 4.66001 V
** VoutMin: 0.150001 V
** VcmMax: 3.35001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.89569e+07 muA
** NormalTransistorNmos: 2.96361e+07 muA
** NormalTransistorNmos: 2.96371e+07 muA
** NormalTransistorNmos: 2.96381e+07 muA
** NormalTransistorNmos: 2.96371e+07 muA
** NormalTransistorPmos: -5.92739e+07 muA
** NormalTransistorPmos: -2.96369e+07 muA
** NormalTransistorPmos: -2.96369e+07 muA
** NormalTransistorNmos: 9.08191e+07 muA
** NormalTransistorPmos: -9.08199e+07 muA
** DiodeTransistorNmos: 1.89561e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.09201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.80401  V


.END