** Name: two_stage_single_output_op_amp_73_7

.MACRO two_stage_single_output_op_amp_73_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=30e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=23e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=22e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=540e-6
m7 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=6e-6 W=57e-6
m8 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
m9 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=31e-6
m11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=31e-6
m12 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=14e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=128e-6
m14 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=180e-6
m15 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=577e-6
m16 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=154e-6
m17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=180e-6
m18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=89e-6
m19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=89e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.20001e-12
.EOM two_stage_single_output_op_amp_73_7

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 8.69601 mW
** Area: 5488 (mu_m)^2
** Transit frequency: 4.34301 MHz
** Transit frequency with error factor: 4.34296 MHz
** Slew rate: 3.88808 V/mu_s
** Phase margin: 60.1606°
** CMRR: 144 dB
** VoutMax: 4.25 V
** VoutMin: 0.170001 V
** VcmMax: 5.13001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorPmos: -2.6638e+08 muA
** NormalTransistorPmos: -7.09669e+07 muA
** NormalTransistorPmos: -2.43679e+07 muA
** NormalTransistorPmos: -4.10879e+07 muA
** NormalTransistorPmos: -2.43679e+07 muA
** NormalTransistorPmos: -4.10879e+07 muA
** NormalTransistorNmos: 2.43671e+07 muA
** NormalTransistorNmos: 2.43671e+07 muA
** DiodeTransistorNmos: 2.43671e+07 muA
** NormalTransistorNmos: 3.34371e+07 muA
** NormalTransistorNmos: 3.34361e+07 muA
** NormalTransistorNmos: 1.67191e+07 muA
** NormalTransistorNmos: 1.67191e+07 muA
** NormalTransistorNmos: 1.29964e+09 muA
** NormalTransistorPmos: -1.29963e+09 muA
** DiodeTransistorNmos: 2.66381e+08 muA
** DiodeTransistorNmos: 7.09661e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.15901  V
** outVoltageBiasXXnXX1: 0.964001  V
** outVoltageBiasXXnXX2: 0.573001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.560001  V
** innerStageBias: 0.391001  V
** out1: 1.13901  V
** sourceGCC1: 4.03801  V
** sourceGCC2: 4.03801  V
** sourceTransconductance: 1.89901  V


.END