.suckt  two_stage_single_output_op_amp_141_2 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m3 FirstStageYinnerLoad1 FirstStageYinnerLoad1 sourceNmos sourceNmos nmos
m4 outFirstStage FirstStageYinnerLoad1 sourceNmos sourceNmos nmos
m5 FirstStageYinnerLoad1 ibias sourcePmos sourcePmos pmos
m6 outFirstStage ibias sourcePmos sourcePmos pmos
m7 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m8 FirstStageYinnerLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c2 out sourceNmos 
m10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m12 out ibias sourcePmos sourcePmos pmos
m13 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m14 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m15 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_141_2

