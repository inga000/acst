** Name: two_stage_single_output_op_amp_60_2

.MACRO two_stage_single_output_op_amp_60_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=97e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=46e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=14e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=542e-6
m7 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=433e-6
m8 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=519e-6
m9 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=519e-6
m10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=235e-6
m11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=600e-6
m12 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=433e-6
m13 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
m14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=46e-6
m15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=52e-6
m16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=52e-6
m17 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=542e-6
m18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
m19 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=74e-6
m20 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=534e-6
m21 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=8e-6 W=332e-6
m22 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=25e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 15.5e-12
.EOM two_stage_single_output_op_amp_60_2

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 6.09701 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 4.83701 MHz
** Transit frequency with error factor: 4.8366 MHz
** Slew rate: 12.6262 V/mu_s
** Phase margin: 60.1606°
** CMRR: 122 dB
** VoutMax: 4.69001 V
** VoutMin: 0.340001 V
** VcmMax: 3.04001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 6.34901e+06 muA
** NormalTransistorPmos: -2.11269e+07 muA
** NormalTransistorPmos: -6.15839e+07 muA
** NormalTransistorNmos: 2.06177e+08 muA
** NormalTransistorNmos: 3.29504e+08 muA
** NormalTransistorNmos: 2.06177e+08 muA
** NormalTransistorNmos: 3.29504e+08 muA
** NormalTransistorPmos: -2.06176e+08 muA
** NormalTransistorPmos: -2.06176e+08 muA
** DiodeTransistorPmos: -2.06176e+08 muA
** NormalTransistorPmos: -2.46656e+08 muA
** DiodeTransistorPmos: -2.46657e+08 muA
** NormalTransistorPmos: -1.23327e+08 muA
** NormalTransistorPmos: -1.23327e+08 muA
** NormalTransistorNmos: 4.51277e+08 muA
** NormalTransistorNmos: 4.51276e+08 muA
** NormalTransistorPmos: -4.51276e+08 muA
** DiodeTransistorNmos: 2.11261e+07 muA
** DiodeTransistorNmos: 6.15831e+07 muA
** DiodeTransistorPmos: -6.34999e+06 muA
** NormalTransistorPmos: -6.35099e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.55201  V
** outSourceVoltageBiasXXpXX1: 4.27601  V
** outVoltageBiasXXnXX1: 0.905001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 3.72501  V
** out1: 2.63201  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.57701  V
** innerTransconductance: 0.311001  V
** inner: 4.27501  V


.END