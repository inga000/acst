** Name: two_stage_single_output_op_amp_50_4

.MACRO two_stage_single_output_op_amp_50_4 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=151e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=55e-6
m3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=173e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=10e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
m6 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=4e-6
m7 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=4e-6
m8 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=76e-6
m9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=245e-6
m10 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=8e-6 W=139e-6
m11 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=151e-6
m12 FirstStageYinnerLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=427e-6
m13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=26e-6
m14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=26e-6
m15 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=185e-6
m16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=119e-6
m17 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=4e-6 W=358e-6
m18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=427e-6
m19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=38e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_50_4

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 5.07101 mW
** Area: 11411 (mu_m)^2
** Transit frequency: 3.38801 MHz
** Transit frequency with error factor: 3.38531 MHz
** Slew rate: 9.30539 V/mu_s
** Phase margin: 61.8795°
** CMRR: 100 dB
** VoutMax: 3.15001 V
** VoutMin: 0.710001 V
** VcmMax: 4.66001 V
** VcmMin: 1.01001 V


** Expected Currents: 
** NormalTransistorPmos: -2.98843e+08 muA
** NormalTransistorPmos: -9.64569e+07 muA
** NormalTransistorPmos: -4.31289e+07 muA
** NormalTransistorPmos: -6.46919e+07 muA
** NormalTransistorPmos: -4.31309e+07 muA
** NormalTransistorPmos: -6.46959e+07 muA
** DiodeTransistorNmos: 4.31301e+07 muA
** NormalTransistorNmos: 4.31301e+07 muA
** NormalTransistorNmos: 4.31271e+07 muA
** NormalTransistorNmos: 2.15641e+07 muA
** NormalTransistorNmos: 2.15641e+07 muA
** NormalTransistorNmos: 4.69596e+08 muA
** NormalTransistorNmos: 4.69595e+08 muA
** NormalTransistorPmos: -4.69595e+08 muA
** NormalTransistorPmos: -4.69594e+08 muA
** DiodeTransistorNmos: 2.98844e+08 muA
** DiodeTransistorNmos: 9.64561e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.64701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11801  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXnXX2: 0.568001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.558001  V
** sourceGCC1: 3.36101  V
** sourceGCC2: 3.36101  V
** sourceTransconductance: 1.65601  V
** innerStageBias: 3.75101  V
** innerTransconductance: 0.150001  V


.END