.suckt  symmetrical_op_amp43 ibias in1 in2 out sourceNmos sourcePmos
m1 outFirstStage outFirstStage sourceNmos sourceNmos nmos
m2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m3 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m5 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m6 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c1 out sourceNmos 
m7 out outFirstStage sourceNmos sourceNmos nmos
m8 out innerComplementarySecondStage sourcePmos sourcePmos pmos
m9 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos
m10 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m11 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m12 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end symmetrical_op_amp43

