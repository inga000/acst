** Name: two_stage_single_output_op_amp_62_10

.MACRO two_stage_single_output_op_amp_62_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=35e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=85e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=417e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=20e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=201e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=91e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=149e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=149e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=509e-6
mFoldedCascodeFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=91e-6
mMainBias12 outVoltageBiasXXpXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=106e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=417e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=138e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=138e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=201e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=389e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mMainBias19 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=364e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=560e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=69e-6
mMainBias22 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=162e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.3001e-12
.EOM two_stage_single_output_op_amp_62_10

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 5.78001 mW
** Area: 13338 (mu_m)^2
** Transit frequency: 3.94401 MHz
** Transit frequency with error factor: 3.94444 MHz
** Slew rate: 6.32499 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 4.52001 V
** VoutMin: 0.150001 V
** VcmMax: 3 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -1.84916e+08 muA
** NormalTransistorPmos: -8.09479e+07 muA
** NormalTransistorNmos: 9.06881e+07 muA
** NormalTransistorNmos: 1.41896e+08 muA
** NormalTransistorNmos: 9.06881e+07 muA
** NormalTransistorNmos: 1.41896e+08 muA
** DiodeTransistorPmos: -9.06889e+07 muA
** NormalTransistorPmos: -9.06889e+07 muA
** NormalTransistorPmos: -9.06889e+07 muA
** NormalTransistorPmos: -1.02411e+08 muA
** DiodeTransistorPmos: -1.0241e+08 muA
** NormalTransistorPmos: -5.12059e+07 muA
** NormalTransistorPmos: -5.12059e+07 muA
** NormalTransistorNmos: 4.84729e+08 muA
** NormalTransistorPmos: -4.84728e+08 muA
** NormalTransistorPmos: -4.84729e+08 muA
** DiodeTransistorNmos: 1.84917e+08 muA
** DiodeTransistorNmos: 8.09471e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 3.28801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.02001  V
** out: 2.5  V
** outFirstStage: 4.17101  V
** outSourceVoltageBiasXXpXX1: 4.14501  V
** outVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.52001  V
** out1: 4.16501  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.35101  V
** innerTransconductance: 4.46901  V
** inner: 4.14101  V


.END