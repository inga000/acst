** Name: symmetrical_op_amp184

.MACRO symmetrical_op_amp184 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias4 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
mSymmetricalFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=238e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=55e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=88e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=150e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=88e-6
mMainBias12 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mSymmetricalFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=33e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=33e-6
mSymmetricalFirstStageLoad18 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=415e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor19 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=528e-6
mSecondStage1Transconductor20 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=528e-6
mSymmetricalFirstStageLoad21 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=415e-6
mMainBias22 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=32e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp184

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 4.68301 mW
** Area: 4035 (mu_m)^2
** Transit frequency: 22.4061 MHz
** Transit frequency with error factor: 22.4063 MHz
** Slew rate: 21.2867 V/mu_s
** Phase margin: 80.7871°
** CMRR: 143 dB
** negPSRR: 118 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 0.680001 V
** VcmMax: 4.81001 V
** VcmMin: 1.65001 V


** Expected Currents: 
** NormalTransistorNmos: 9.91101e+06 muA
** NormalTransistorNmos: 9.95231e+07 muA
** NormalTransistorPmos: -5.31659e+07 muA
** NormalTransistorPmos: -1.67608e+08 muA
** NormalTransistorPmos: -1.67609e+08 muA
** NormalTransistorPmos: -1.67608e+08 muA
** NormalTransistorPmos: -1.67609e+08 muA
** NormalTransistorNmos: 3.35216e+08 muA
** NormalTransistorNmos: 3.35215e+08 muA
** NormalTransistorNmos: 1.67609e+08 muA
** NormalTransistorNmos: 1.67609e+08 muA
** NormalTransistorNmos: 2.14439e+08 muA
** NormalTransistorNmos: 2.14438e+08 muA
** NormalTransistorPmos: -2.14438e+08 muA
** NormalTransistorPmos: -2.14438e+08 muA
** DiodeTransistorNmos: 2.14439e+08 muA
** NormalTransistorPmos: -2.14438e+08 muA
** NormalTransistorPmos: -2.14438e+08 muA
** DiodeTransistorNmos: 5.31651e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.91199e+06 muA
** DiodeTransistorPmos: -9.95239e+07 muA


** Expected Voltages: 
** ibias: 0.629001  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.863001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 1.09201  V
** outVoltageBiasXXpXX0: 3.68801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.224001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.461001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END