** Name: two_stage_single_output_op_amp_71_4

.MACRO two_stage_single_output_op_amp_71_4 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=13e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=50e-6
m3 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=193e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=19e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m6 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=556e-6
m7 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=193e-6
m8 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=310e-6
m9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=29e-6
m10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=29e-6
m11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=587e-6
m12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=370e-6
m13 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=597e-6
m14 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=413e-6
m15 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
m16 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=48e-6
m17 FirstStageYinnerLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=413e-6
m18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=365e-6
m19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=365e-6
m20 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=542e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 20.3001e-12
.EOM two_stage_single_output_op_amp_71_4

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 7.10501 mW
** Area: 14350 (mu_m)^2
** Transit frequency: 3.36501 MHz
** Transit frequency with error factor: 3.35516 MHz
** Slew rate: 10.6664 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 3.97001 V
** VoutMin: 0.540001 V
** VcmMax: 5.17001 V
** VcmMin: 1.84001 V


** Expected Currents: 
** NormalTransistorPmos: -6.26059e+07 muA
** NormalTransistorPmos: -4.86659e+07 muA
** NormalTransistorPmos: -2.17986e+08 muA
** NormalTransistorPmos: -3.70064e+08 muA
** NormalTransistorPmos: -2.17986e+08 muA
** NormalTransistorPmos: -3.70064e+08 muA
** DiodeTransistorNmos: 2.17987e+08 muA
** NormalTransistorNmos: 2.17987e+08 muA
** NormalTransistorNmos: 3.04154e+08 muA
** NormalTransistorNmos: 3.04153e+08 muA
** NormalTransistorNmos: 1.52078e+08 muA
** NormalTransistorNmos: 1.52078e+08 muA
** NormalTransistorNmos: 5.49523e+08 muA
** NormalTransistorNmos: 5.49522e+08 muA
** NormalTransistorPmos: -5.49522e+08 muA
** NormalTransistorPmos: -5.49521e+08 muA
** DiodeTransistorNmos: 6.26051e+07 muA
** DiodeTransistorNmos: 4.86651e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.46301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.700001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.941001  V
** outVoltageBiasXXnXX2: 0.557001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.710001  V
** innerStageBias: 0.361001  V
** sourceGCC1: 4.19801  V
** sourceGCC2: 4.19801  V
** sourceTransconductance: 1.38801  V
** innerStageBias: 4.25301  V
** innerTransconductance: 0.295001  V


.END