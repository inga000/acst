** Name: two_stage_single_output_op_amp_82_9

.MACRO two_stage_single_output_op_amp_82_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=24e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=24e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=74e-6
mMainBias4 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=6e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=240e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=24e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=16e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=12e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=74e-6
mMainBias14 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=10e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=240e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=43e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=78e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=78e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=472e-6
mFoldedCascodeFirstStageLoad21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=43e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=395e-6
mMainBias23 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.5e-12
.EOM two_stage_single_output_op_amp_82_9

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 11.1581 mW
** Area: 5823 (mu_m)^2
** Transit frequency: 6.38601 MHz
** Transit frequency with error factor: 6.38575 MHz
** Slew rate: 4.39361 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 4.25 V
** VoutMin: 1.77001 V
** VcmMax: 5.17001 V
** VcmMin: 1.47001 V


** Expected Currents: 
** NormalTransistorPmos: -4.00481e+08 muA
** NormalTransistorPmos: -6.59019e+07 muA
** NormalTransistorPmos: -4.62099e+07 muA
** NormalTransistorPmos: -7.90819e+07 muA
** NormalTransistorPmos: -4.62099e+07 muA
** NormalTransistorPmos: -7.90819e+07 muA
** DiodeTransistorNmos: 4.62091e+07 muA
** NormalTransistorNmos: 4.62081e+07 muA
** NormalTransistorNmos: 4.62091e+07 muA
** DiodeTransistorNmos: 4.62081e+07 muA
** NormalTransistorNmos: 6.57411e+07 muA
** DiodeTransistorNmos: 6.57401e+07 muA
** NormalTransistorNmos: 3.28711e+07 muA
** NormalTransistorNmos: 3.28711e+07 muA
** NormalTransistorNmos: 1.58699e+09 muA
** DiodeTransistorNmos: 1.58699e+09 muA
** NormalTransistorPmos: -1.58698e+09 muA
** DiodeTransistorNmos: 4.00482e+08 muA
** NormalTransistorNmos: 4.00481e+08 muA
** DiodeTransistorNmos: 6.59011e+07 muA
** NormalTransistorNmos: 6.59001e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.31801  V
** outInputVoltageBiasXXnXX2: 2.17401  V
** outSourceVoltageBiasXXnXX1: 0.659001  V
** outSourceVoltageBiasXXnXX2: 1.08701  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.856001  V
** innerTransistorStack2Load2: 0.856001  V
** out1: 1.41201  V
** sourceGCC1: 4.21701  V
** sourceGCC2: 4.21701  V
** sourceTransconductance: 1.93901  V
** inner: 0.659001  V
** inner: 1.08301  V


.END