** Name: two_stage_single_output_op_amp_19_1

.MACRO two_stage_single_output_op_amp_19_1 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=12e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=49e-6
m3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
m5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=35e-6
m6 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=153e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=320e-6
m8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=10e-6 W=120e-6
m9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
m10 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
m11 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=203e-6
m12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=45e-6
m13 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
m14 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=45e-6
m15 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=91e-6
m16 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=167e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 5.20001e-12
.EOM two_stage_single_output_op_amp_19_1

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 1.12401 mW
** Area: 6341 (mu_m)^2
** Transit frequency: 3.10301 MHz
** Transit frequency with error factor: 3.09609 MHz
** Slew rate: 4.01367 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** negPSRR: 99 dB
** posPSRR: 205 dB
** VoutMax: 4.83001 V
** VoutMin: 0.150001 V
** VcmMax: 3.09001 V
** VcmMin: 0.140001 V


** Expected Currents: 
** NormalTransistorNmos: 3.66101e+07 muA
** NormalTransistorPmos: -1.17169e+07 muA
** NormalTransistorPmos: -9.16999e+06 muA
** DiodeTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28571e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorPmos: -4.57129e+07 muA
** NormalTransistorPmos: -4.57139e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorNmos: 1.01582e+08 muA
** NormalTransistorPmos: -1.01581e+08 muA
** DiodeTransistorNmos: 1.17161e+07 muA
** DiodeTransistorNmos: 9.16901e+06 muA
** DiodeTransistorPmos: -3.66109e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXpXX1: 4.09301  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerStageBias: 4.83201  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.50801  V


.END