** Name: two_stage_single_output_op_amp_50_8

.MACRO two_stage_single_output_op_amp_50_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=18e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=23e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=24e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageTransconductor6 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=60e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=60e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=565e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=550e-6
mFoldedCascodeFirstStageLoad11 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=18e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=295e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=134e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=134e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=231e-6
mFoldedCascodeFirstStageLoad16 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=295e-6
mMainBias17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=181e-6
mMainBias18 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=99e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.5e-12
.EOM two_stage_single_output_op_amp_50_8

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 7.28601 mW
** Area: 7295 (mu_m)^2
** Transit frequency: 3.39201 MHz
** Transit frequency with error factor: 3.3885 MHz
** Slew rate: 3.76925 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.25 V
** VoutMin: 0.380001 V
** VcmMax: 5.12001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorPmos: -8.68879e+07 muA
** NormalTransistorPmos: -4.75169e+07 muA
** NormalTransistorPmos: -3.99359e+07 muA
** NormalTransistorPmos: -6.50289e+07 muA
** NormalTransistorPmos: -3.99359e+07 muA
** NormalTransistorPmos: -6.50289e+07 muA
** DiodeTransistorNmos: 3.99351e+07 muA
** NormalTransistorNmos: 3.99351e+07 muA
** NormalTransistorNmos: 5.01831e+07 muA
** NormalTransistorNmos: 2.50921e+07 muA
** NormalTransistorNmos: 2.50921e+07 muA
** NormalTransistorNmos: 1.17272e+09 muA
** NormalTransistorNmos: 1.17272e+09 muA
** NormalTransistorPmos: -1.17271e+09 muA
** DiodeTransistorNmos: 8.68871e+07 muA
** DiodeTransistorNmos: 4.75161e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** outVoltageBiasXXnXX1: 0.987001  V
** outVoltageBiasXXnXX2: 0.562001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.915001  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.87201  V
** innerStageBias: 0.357001  V


.END