** Name: symmetrical_op_amp147

.MACRO symmetrical_op_amp147 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
m2 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=1e-6 W=235e-6
m3 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=235e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m6 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=125e-6
m7 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=1e-6 W=132e-6
m8 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=132e-6
m9 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=125e-6
m10 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=475e-6
m11 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=476e-6
m12 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=545e-6
m13 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=545e-6
m14 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=516e-6
m15 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=235e-6
m16 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=516e-6
m17 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=161e-6
m18 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
m19 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=551e-6
m20 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=235e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp147

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 7.43501 mW
** Area: 13056 (mu_m)^2
** Transit frequency: 15.2291 MHz
** Transit frequency with error factor: 15.2287 MHz
** Slew rate: 34.4601 V/mu_s
** Phase margin: 69.328°
** CMRR: 143 dB
** negPSRR: 46 dB
** posPSRR: 73 dB
** VoutMax: 3.86001 V
** VoutMin: 0.330001 V
** VcmMax: 3.03001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.63233e+08 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04163e+08 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04163e+08 muA
** NormalTransistorPmos: -6.08327e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorNmos: 3.46009e+08 muA
** NormalTransistorNmos: 3.46008e+08 muA
** NormalTransistorPmos: -3.46008e+08 muA
** DiodeTransistorPmos: -3.46009e+08 muA
** DiodeTransistorPmos: -3.49502e+08 muA
** NormalTransistorPmos: -3.49503e+08 muA
** NormalTransistorNmos: 3.49503e+08 muA
** NormalTransistorNmos: 3.49502e+08 muA
** DiodeTransistorNmos: 1.63234e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 4.14801  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 3.29601  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.731001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.22101  V
** innerTransistorStack1Load1: 0.156001  V
** innerTransistorStack2Load1: 0.156001  V
** sourceTransconductance: 3.42601  V
** innerTransconductance: 0.150001  V
** inner: 4.14801  V
** inner: 0.150001  V


.END