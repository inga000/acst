.suckt  one_stage_single_output_op_amp97 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mMainBias2 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mTelescopicFirstStageLoad3 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mTelescopicFirstStageLoad4 out outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos
mTelescopicFirstStageLoad7 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos
mTelescopicFirstStageLoad8 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos
mTelescopicFirstStageStageBias9 sourceTransconductance ibias sourceNmos sourceNmos nmos
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
cLoadCapacitor1 out sourceNmos 
mMainBias12 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
mMainBias13 ibias ibias sourceNmos sourceNmos nmos
mMainBias14 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end one_stage_single_output_op_amp97

