.suckt  two_stage_single_output_op_amp_127_7 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 FirstStageYinnerLoad1 FirstStageYinnerLoad1 sourcePmos sourcePmos pmos
m3 outFirstStage FirstStageYinnerLoad1 sourcePmos sourcePmos pmos
m4 FirstStageYinnerLoad1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m5 outFirstStage outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m6 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m7 FirstStageYinnerLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c2 out sourceNmos 
m9 out outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m10 out outFirstStage sourcePmos sourcePmos pmos
m11 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m12 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_127_7

