.suckt  two_stage_fully_differential_op_amp_43_6 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 outInputVoltageBiasXXpXX3 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m4 outVoltageBiasXXpXX4 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m5 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m6 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m7 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m8 outFeedback outFeedback sourceNmos sourceNmos nmos
m9 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m10 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m11 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m15 out1FirstStage outVoltageBiasXXpXX4 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m16 out2FirstStage outVoltageBiasXXpXX4 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m17 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m18 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m19 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m20 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m21 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m22 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m23 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m24 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m25 out1 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m26 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m27 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m28 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m29 out2 outInputVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos
m30 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m31 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m32 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m33 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m34 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m35 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m36 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m37 outInputVoltageBiasXXpXX3 outInputVoltageBiasXXpXX3 VoltageBiasXXpXX3Yinner VoltageBiasXXpXX3Yinner pmos
m38 VoltageBiasXXpXX3Yinner outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m39 outVoltageBiasXXpXX4 outVoltageBiasXXpXX4 sourceTransconductance sourceTransconductance pmos
m40 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_43_6

