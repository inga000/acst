.suckt  two_stage_single_output_op_amp_31_7 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_3 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_4 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_StageBias_6 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_SingleOutput_FirstStage_StageBias_7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Transconductor_8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_SingleOutput_FirstStage_Transconductor_9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_StageBias_10 out ibias sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_Transconductor_11 out outFirstStage sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_12 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_13 ibias ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_14 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_31_7

