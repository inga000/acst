** Name: two_stage_single_output_op_amp_196_8

.MACRO two_stage_single_output_op_amp_196_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=7e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=11e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=6e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=68e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mMainBias7 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=91e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=19e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=68e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=598e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=6e-6
mSecondStage1StageBias13 out inputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=7e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=19e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=563e-6
mMainBias17 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=189e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=230e-6
mSimpleFirstStageLoad19 outFirstStage ibias sourcePmos sourcePmos pmos4 L=4e-6 W=563e-6
mMainBias20 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=29e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.60001e-12
.EOM two_stage_single_output_op_amp_196_8

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 6.56401 mW
** Area: 8392 (mu_m)^2
** Transit frequency: 4.39301 MHz
** Transit frequency with error factor: 4.38268 MHz
** Slew rate: 4.14033 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 0.700001 V
** VcmMax: 5.25 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorPmos: -3.21599e+06 muA
** NormalTransistorPmos: -2.09519e+07 muA
** DiodeTransistorNmos: 4.33721e+07 muA
** DiodeTransistorNmos: 4.33711e+07 muA
** NormalTransistorNmos: 4.33701e+07 muA
** NormalTransistorNmos: 4.33711e+07 muA
** NormalTransistorPmos: -6.14649e+07 muA
** NormalTransistorPmos: -6.14649e+07 muA
** NormalTransistorNmos: 3.61871e+07 muA
** DiodeTransistorNmos: 3.61861e+07 muA
** NormalTransistorNmos: 1.80941e+07 muA
** NormalTransistorNmos: 1.80941e+07 muA
** NormalTransistorNmos: 1.1457e+09 muA
** NormalTransistorNmos: 1.1457e+09 muA
** NormalTransistorPmos: -1.14569e+09 muA
** DiodeTransistorNmos: 3.21501e+06 muA
** NormalTransistorNmos: 3.21401e+06 muA
** DiodeTransistorNmos: 2.09511e+07 muA
** DiodeTransistorNmos: 2.09511e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.11001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.16401  V
** outSourceVoltageBiasXXnXX1: 0.582001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.12401  V
** innerTransistorStack2Load1: 1.125  V
** out1: 2.19501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.555001  V
** inner: 0.581001  V


.END