** Name: two_stage_single_output_op_amp_9_11

.MACRO two_stage_single_output_op_amp_9_11 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=94e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=468e-6
mMainBias4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1StageBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=119e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=65e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
mMainBias9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=37e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=8e-6 W=557e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=119e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=50e-6
mSimpleFirstStageLoad13 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=468e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=395e-6
mSecondStage1Transconductor15 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=199e-6
mMainBias17 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=59e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16e-12
.EOM two_stage_single_output_op_amp_9_11

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 9.80401 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 7.10901 MHz
** Transit frequency with error factor: 7.10524 MHz
** Slew rate: 7.96996 V/mu_s
** Phase margin: 60.1606°
** CMRR: 106 dB
** negPSRR: 110 dB
** posPSRR: 100 dB
** VoutMax: 4.25 V
** VoutMin: 0.670001 V
** VcmMax: 4.44001 V
** VcmMin: 0.800001 V


** Expected Currents: 
** NormalTransistorNmos: 7.44871e+07 muA
** NormalTransistorNmos: 1.00659e+08 muA
** NormalTransistorPmos: -4.39437e+08 muA
** NormalTransistorPmos: -6.41339e+07 muA
** NormalTransistorPmos: -6.41339e+07 muA
** DiodeTransistorPmos: -6.41339e+07 muA
** NormalTransistorNmos: 1.28267e+08 muA
** NormalTransistorNmos: 6.41331e+07 muA
** NormalTransistorNmos: 6.41331e+07 muA
** NormalTransistorNmos: 1.20791e+09 muA
** NormalTransistorNmos: 1.20791e+09 muA
** NormalTransistorPmos: -1.2079e+09 muA
** NormalTransistorPmos: -1.2079e+09 muA
** DiodeTransistorNmos: 4.39438e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -7.44879e+07 muA
** DiodeTransistorPmos: -1.00658e+08 muA


** Expected Voltages: 
** ibias: 0.622001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.78801  V
** out: 2.5  V
** outFirstStage: 4.02101  V
** outVoltageBiasXXnXX1: 1.07301  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.22101  V
** out1: 3.46701  V
** sourceTransconductance: 1.91601  V
** innerStageBias: 0.217001  V
** innerTransconductance: 4.58501  V


.END