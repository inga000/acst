** Name: two_stage_single_output_op_amp_13_8

.MACRO two_stage_single_output_op_amp_13_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=59e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=59e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=27e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=8e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=170e-6
mMainBias9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=196e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=8e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=59e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=334e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=59e-6
mMainBias15 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=100e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_13_8

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 2.53701 mW
** Area: 6781 (mu_m)^2
** Transit frequency: 2.54301 MHz
** Transit frequency with error factor: 2.53915 MHz
** Slew rate: 5.96466 V/mu_s
** Phase margin: 61.8795°
** CMRR: 100 dB
** negPSRR: 90 dB
** posPSRR: 86 dB
** VoutMax: 4.25 V
** VoutMin: 0.660001 V
** VcmMax: 3.76001 V
** VcmMin: 1.12001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00011e+07 muA
** NormalTransistorPmos: -3.66209e+07 muA
** DiodeTransistorPmos: -1.34799e+07 muA
** NormalTransistorPmos: -1.34809e+07 muA
** NormalTransistorPmos: -1.34799e+07 muA
** DiodeTransistorPmos: -1.34809e+07 muA
** NormalTransistorNmos: 2.69591e+07 muA
** NormalTransistorNmos: 1.34791e+07 muA
** NormalTransistorNmos: 1.34791e+07 muA
** NormalTransistorNmos: 4.23904e+08 muA
** NormalTransistorNmos: 4.23903e+08 muA
** NormalTransistorPmos: -4.23903e+08 muA
** DiodeTransistorNmos: 3.66201e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.00019e+07 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.00501  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 1.06601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.11501  V
** innerTransistorStack1Load1: 4.11401  V
** out1: 3.35501  V
** sourceTransconductance: 1.72001  V
** innerStageBias: 0.342001  V


.END