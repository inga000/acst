** Name: one_stage_single_output_op_amp47

.MACRO one_stage_single_output_op_amp47 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=13e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=113e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=449e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=449e-6
mMainBias8 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=66e-6
mMainBias9 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=22e-6
mFoldedCascodeFirstStageLoad10 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=113e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=292e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=126e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=126e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=126e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=126e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=54e-6
mFoldedCascodeFirstStageLoad17 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=292e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp47

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 1.93001 mW
** Area: 8363 (mu_m)^2
** Transit frequency: 5.69301 MHz
** Transit frequency with error factor: 5.6935 MHz
** Slew rate: 5.65981 V/mu_s
** Phase margin: 84.2249°
** CMRR: 138 dB
** VoutMax: 4.47001 V
** VoutMin: 0.800001 V
** VcmMax: 3.68001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.53821e+07 muA
** NormalTransistorNmos: 8.46401e+06 muA
** NormalTransistorNmos: 1.13698e+08 muA
** NormalTransistorNmos: 1.71037e+08 muA
** NormalTransistorNmos: 1.13698e+08 muA
** NormalTransistorNmos: 1.71037e+08 muA
** NormalTransistorPmos: -1.13697e+08 muA
** NormalTransistorPmos: -1.13698e+08 muA
** NormalTransistorPmos: -1.13697e+08 muA
** NormalTransistorPmos: -1.13698e+08 muA
** NormalTransistorPmos: -1.1468e+08 muA
** NormalTransistorPmos: -5.73399e+07 muA
** NormalTransistorPmos: -5.73399e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.53829e+07 muA
** DiodeTransistorPmos: -8.46499e+06 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** inputVoltageBiasXXpXX2: 3.83701  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.11701  V
** innerTransistorStack1Load2: 4.45801  V
** innerTransistorStack2Load2: 4.45801  V
** sourceGCC1: 0.523001  V
** sourceGCC2: 0.523001  V
** sourceTransconductance: 3.22301  V


.END