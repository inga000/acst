** Name: two_stage_single_output_op_amp_109_1

.MACRO two_stage_single_output_op_amp_109_1 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=419e-6
m2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=58e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=58e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
m5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=79e-6
m6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=52e-6
m7 inputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=565e-6
m8 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=150e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=3e-6 W=58e-6
m10 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=421e-6
m11 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=58e-6
m12 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=599e-6
m13 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=41e-6
m14 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=479e-6
m15 sourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=427e-6
m16 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
m17 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=41e-6
m18 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=20e-6
m19 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=20e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.80001e-12
.EOM two_stage_single_output_op_amp_109_1

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 7.39101 mW
** Area: 14934 (mu_m)^2
** Transit frequency: 5.34001 MHz
** Transit frequency with error factor: 5.34014 MHz
** Slew rate: 15.1174 V/mu_s
** Phase margin: 60.1606°
** CMRR: 127 dB
** VoutMax: 4.81001 V
** VoutMin: 0.300001 V
** VcmMax: 3.01001 V
** VcmMin: 0.860001 V


** Expected Currents: 
** NormalTransistorNmos: 3.05076e+08 muA
** NormalTransistorNmos: 4.03224e+08 muA
** NormalTransistorPmos: -2.99028e+08 muA
** NormalTransistorPmos: -3.68239e+07 muA
** NormalTransistorPmos: -3.68239e+07 muA
** DiodeTransistorNmos: 3.68231e+07 muA
** NormalTransistorNmos: 3.68231e+07 muA
** NormalTransistorNmos: 3.68231e+07 muA
** DiodeTransistorNmos: 3.68231e+07 muA
** NormalTransistorPmos: -3.78724e+08 muA
** NormalTransistorPmos: -3.78723e+08 muA
** NormalTransistorPmos: -3.68249e+07 muA
** NormalTransistorPmos: -3.68249e+07 muA
** NormalTransistorNmos: 3.77155e+08 muA
** NormalTransistorPmos: -3.77154e+08 muA
** DiodeTransistorNmos: 2.99029e+08 muA
** DiodeTransistorPmos: -3.05075e+08 muA
** DiodeTransistorPmos: -4.03223e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.89901  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outVoltageBiasXXnXX0: 0.666001  V
** outVoltageBiasXXpXX1: 2.13801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.51601  V
** innerSourceLoad2: 0.555001  V
** innerStageBias: 4.68501  V
** innerTransistorStack1Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 3.01801  V
** sourceGCC2: 3.01801  V


.END