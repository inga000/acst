.suckt  symmetrical_op_amp1 ibias in1 in2 out sourceNmos sourcePmos
mSymmetricalFirstStageLoad1 outFirstStage outFirstStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageLoad2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageStageBias3 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSymmetricalFirstStageTransconductor4 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSymmetricalFirstStageTransconductor5 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias7 out innerComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias8 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mMainBias10 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp1

