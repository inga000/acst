** Name: two_stage_single_output_op_amp_3_5

.MACRO two_stage_single_output_op_amp_3_5 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=30e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=9e-6 W=192e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=6e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=204e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=30e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=192e-6
mSimpleFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=14e-6
mMainBias10 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=20e-6
mSimpleFirstStageTransconductor11 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=23e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=9e-6 W=369e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=6e-6
mMainBias14 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=9e-6 W=248e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=204e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=23e-6
mMainBias17 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=9e-6 W=47e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_3_5

** Expected Performance Values: 
** Gain: 108 dB
** Power consumption: 1.21401 mW
** Area: 10912 (mu_m)^2
** Transit frequency: 4.41601 MHz
** Transit frequency with error factor: 4.4134 MHz
** Slew rate: 4.22426 V/mu_s
** Phase margin: 67.0361°
** CMRR: 106 dB
** negPSRR: 108 dB
** posPSRR: 222 dB
** VoutMax: 3.43001 V
** VoutMin: 0.150001 V
** VcmMax: 4.12001 V
** VcmMin: 0.150001 V


** Expected Currents: 
** NormalTransistorNmos: 5.44701e+06 muA
** NormalTransistorPmos: -2.47299e+06 muA
** NormalTransistorPmos: -1.29959e+07 muA
** DiodeTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorPmos: -1.90509e+07 muA
** NormalTransistorPmos: -9.52499e+06 muA
** NormalTransistorPmos: -9.52499e+06 muA
** NormalTransistorNmos: 1.82918e+08 muA
** NormalTransistorPmos: -1.82917e+08 muA
** DiodeTransistorPmos: -1.82918e+08 muA
** DiodeTransistorNmos: 2.47201e+06 muA
** DiodeTransistorNmos: 1.29951e+07 muA
** DiodeTransistorPmos: -5.44799e+06 muA
** NormalTransistorPmos: -5.44899e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.710001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.86601  V
** outSourceVoltageBiasXXpXX1: 3.93301  V
** outVoltageBiasXXnXX0: 0.576001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.21601  V
** inner: 3.93201  V


.END