** Name: symmetrical_op_amp153

.MACRO symmetrical_op_amp153 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=46e-6
mMainBias2 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=20e-6
mSecondStage1StageBias3 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=214e-6
mSymmetricalFirstStageStageBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=63e-6
mSymmetricalFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=42e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=42e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=110e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=110e-6
mSymmetricalFirstStageLoad9 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=44e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=46e-6
mSecondStage1Transconductor11 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=46e-6
mSymmetricalFirstStageLoad12 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=44e-6
mSymmetricalFirstStageStageBias13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=63e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mSymmetricalFirstStageTransconductor15 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=119e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias16 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=214e-6
mSecondStage1StageBias17 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=2e-6 W=153e-6
mSymmetricalFirstStageTransconductor18 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=119e-6
mMainBias19 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=211e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp153

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 1.21201 mW
** Area: 7643 (mu_m)^2
** Transit frequency: 3.43601 MHz
** Transit frequency with error factor: 3.43636 MHz
** Slew rate: 4.18102 V/mu_s
** Phase margin: 66.4632°
** CMRR: 150 dB
** negPSRR: 48 dB
** posPSRR: 55 dB
** VoutMax: 4.03001 V
** VoutMin: 0.400001 V
** VcmMax: 3.09001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.06465e+08 muA
** NormalTransistorNmos: 1.60491e+07 muA
** NormalTransistorNmos: 1.60481e+07 muA
** NormalTransistorNmos: 1.60491e+07 muA
** NormalTransistorNmos: 1.60481e+07 muA
** NormalTransistorPmos: -3.20999e+07 muA
** DiodeTransistorPmos: -3.20989e+07 muA
** NormalTransistorPmos: -1.60499e+07 muA
** NormalTransistorPmos: -1.60499e+07 muA
** NormalTransistorNmos: 4.19011e+07 muA
** NormalTransistorNmos: 4.19021e+07 muA
** NormalTransistorPmos: -4.19019e+07 muA
** DiodeTransistorPmos: -4.19029e+07 muA
** NormalTransistorPmos: -4.19019e+07 muA
** NormalTransistorNmos: 4.19011e+07 muA
** NormalTransistorNmos: 4.19021e+07 muA
** DiodeTransistorNmos: 1.06466e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.28801  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** inStageBiasComplementarySecondStage: 4.20101  V
** innerComplementarySecondStage: 3.46201  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.808001  V
** outSourceVoltageBiasXXpXX1: 4.14501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.242001  V
** innerTransistorStack2Load1: 0.242001  V
** sourceTransconductance: 3.25801  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V
** inner: 4.14101  V


.END