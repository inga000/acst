** Name: two_stage_single_output_op_amp_81_9

.MACRO two_stage_single_output_op_amp_81_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=16e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=16e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=11e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=10e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=534e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=132e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=9e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=28e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=62e-6
mFoldedCascodeFirstStageLoad10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=11e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=11e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=6e-6 W=7e-6
mMainBias14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=10e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=534e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=16e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=147e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=130e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=130e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=196e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=502e-6
mFoldedCascodeFirstStageLoad22 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=147e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=33e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_81_9

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 4.15601 mW
** Area: 14998 (mu_m)^2
** Transit frequency: 2.90101 MHz
** Transit frequency with error factor: 2.90072 MHz
** Slew rate: 6.56198 V/mu_s
** Phase margin: 64.7443°
** CMRR: 137 dB
** VoutMax: 4.25 V
** VoutMin: 1.03001 V
** VcmMax: 5.21001 V
** VcmMin: 1.99001 V


** Expected Currents: 
** NormalTransistorPmos: -1.17299e+07 muA
** NormalTransistorPmos: -6.93979e+07 muA
** NormalTransistorPmos: -2.98509e+07 muA
** NormalTransistorPmos: -4.64629e+07 muA
** NormalTransistorPmos: -2.98509e+07 muA
** NormalTransistorPmos: -4.64629e+07 muA
** DiodeTransistorNmos: 2.98501e+07 muA
** NormalTransistorNmos: 2.98491e+07 muA
** NormalTransistorNmos: 2.98501e+07 muA
** DiodeTransistorNmos: 2.98491e+07 muA
** NormalTransistorNmos: 3.32211e+07 muA
** NormalTransistorNmos: 3.32201e+07 muA
** NormalTransistorNmos: 1.66111e+07 muA
** NormalTransistorNmos: 1.66111e+07 muA
** NormalTransistorNmos: 6.37126e+08 muA
** DiodeTransistorNmos: 6.37125e+08 muA
** NormalTransistorPmos: -6.37125e+08 muA
** DiodeTransistorNmos: 1.17291e+07 muA
** NormalTransistorNmos: 1.17301e+07 muA
** DiodeTransistorNmos: 6.93971e+07 muA
** DiodeTransistorNmos: 6.93961e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.67001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.43601  V
** outSourceVoltageBiasXXnXX1: 0.718001  V
** outSourceVoltageBiasXXnXX2: 0.599001  V
** outSourceVoltageBiasXXpXX1: 4.23701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.683001  V
** innerTransistorStack1Load2: 0.766001  V
** innerTransistorStack2Load2: 0.767001  V
** out1: 1.38101  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.69301  V
** inner: 0.719001  V


.END