** Name: symmetrical_op_amp153

.MACRO symmetrical_op_amp153 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m2 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=33e-6
m3 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=382e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=200e-6
m5 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=2e-6 W=49e-6
m6 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=32e-6
m7 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=49e-6
m8 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=32e-6
m9 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=80e-6
m10 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=80e-6
m11 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=143e-6
m12 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=143e-6
m13 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=382e-6
m14 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=18e-6
m15 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=6e-6 W=159e-6
m16 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=18e-6
m17 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=69e-6
m18 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=200e-6
m19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=33e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp153

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 1.05601 mW
** Area: 11042 (mu_m)^2
** Transit frequency: 2.82201 MHz
** Transit frequency with error factor: 2.82246 MHz
** Slew rate: 5.43482 V/mu_s
** Phase margin: 77.9223°
** CMRR: 144 dB
** negPSRR: 48 dB
** posPSRR: 69 dB
** VoutMax: 3.86001 V
** VoutMin: 0.310001 V
** VcmMax: 3.04001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.08089e+07 muA
** NormalTransistorNmos: 3.07401e+07 muA
** NormalTransistorNmos: 3.07391e+07 muA
** NormalTransistorNmos: 3.07401e+07 muA
** NormalTransistorNmos: 3.07391e+07 muA
** NormalTransistorPmos: -6.14809e+07 muA
** DiodeTransistorPmos: -6.14799e+07 muA
** NormalTransistorPmos: -3.07409e+07 muA
** NormalTransistorPmos: -3.07409e+07 muA
** NormalTransistorNmos: 5.44721e+07 muA
** NormalTransistorNmos: 5.44731e+07 muA
** NormalTransistorPmos: -5.44729e+07 muA
** DiodeTransistorPmos: -5.44739e+07 muA
** NormalTransistorPmos: -5.44749e+07 muA
** NormalTransistorNmos: 5.44741e+07 muA
** NormalTransistorNmos: 5.44731e+07 muA
** DiodeTransistorNmos: 2.08081e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.34801  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** inStageBiasComplementarySecondStage: 4.19901  V
** innerComplementarySecondStage: 3.29501  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.717001  V
** outSourceVoltageBiasXXpXX1: 4.17501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.161001  V
** innerTransistorStack2Load1: 0.161001  V
** sourceTransconductance: 3.37201  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V
** inner: 4.17201  V


.END