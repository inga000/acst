** Name: two_stage_single_output_op_amp_65_9

.MACRO two_stage_single_output_op_amp_65_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=12e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=120e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=9e-6 W=194e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=120e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
mMainBias13 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=32e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=9e-6 W=449e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=42e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=42e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=51e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=48e-6
mFoldedCascodeFirstStageTransconductor19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=48e-6
mFoldedCascodeFirstStageStageBias20 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=52e-6
mMainBias21 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=9e-6 W=445e-6
mSecondStage1Transconductor22 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=467e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=51e-6
mMainBias24 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=9e-6 W=393e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_65_9

** Expected Performance Values: 
** Gain: 135 dB
** Power consumption: 2.21201 mW
** Area: 14994 (mu_m)^2
** Transit frequency: 2.85301 MHz
** Transit frequency with error factor: 2.85275 MHz
** Slew rate: 5.05082 V/mu_s
** Phase margin: 76.7764°
** CMRR: 141 dB
** VoutMax: 4.83001 V
** VoutMin: 0.720001 V
** VcmMax: 3.27001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 6.15631e+07 muA
** NormalTransistorPmos: -2.03989e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorNmos: 2.28181e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 2.28181e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorPmos: -2.28189e+07 muA
** NormalTransistorPmos: -2.28199e+07 muA
** NormalTransistorPmos: -2.28189e+07 muA
** NormalTransistorPmos: -2.28199e+07 muA
** NormalTransistorPmos: -2.29349e+07 muA
** NormalTransistorPmos: -2.29359e+07 muA
** NormalTransistorPmos: -1.14669e+07 muA
** NormalTransistorPmos: -1.14669e+07 muA
** NormalTransistorNmos: 2.49044e+08 muA
** DiodeTransistorNmos: 2.49043e+08 muA
** NormalTransistorPmos: -2.49043e+08 muA
** DiodeTransistorNmos: 2.03981e+07 muA
** NormalTransistorNmos: 2.03971e+07 muA
** DiodeTransistorNmos: 2.28561e+07 muA
** DiodeTransistorNmos: 2.28561e+07 muA
** DiodeTransistorPmos: -6.15639e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.11001  V
** out: 2.5  V
** outFirstStage: 4.26301  V
** outInputVoltageBiasXXnXX1: 1.12201  V
** outSourceVoltageBiasXXnXX1: 0.561001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.89901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.62001  V
** innerTransistorStack1Load2: 4.62101  V
** innerTransistorStack2Load2: 4.62101  V
** out1: 4.26101  V
** sourceGCC1: 0.540001  V
** sourceGCC2: 0.540001  V
** sourceTransconductance: 3.34601  V
** inner: 0.561001  V


.END