.suckt  two_stage_fully_differential_op_amp_53_8 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_3 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_4 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_5 outFeedback outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_6 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackStage_Transconductor_8 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_9 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_10 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FeedbackStage_Transconductor_11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FirstStage_Load_12 out1FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m_FullyDifferential_FirstStage_Load_13 FirstStageYinnerTransistorStack1Load1 outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_14 out2FirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_FullyDifferential_FirstStage_Load_15 FirstStageYinnerTransistorStack2Load1 outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_StageBias_16 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_FullyDifferential_FirstStage_StageBias_17 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Transconductor_18 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_FullyDifferential_FirstStage_Transconductor_19 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_StageBias_20 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias nmos
m_FullyDifferential_SecondStage1_StageBias_21 SecondStage1YinnerStageBias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_Transconductor_22 out1 out1FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_StageBias_23 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias nmos
m_FullyDifferential_SecondStage2_StageBias_24 SecondStage2YinnerStageBias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_Transconductor_25 out2 out2FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_26 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_27 ibias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_28 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_29 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_53_8

