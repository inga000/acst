.suckt  symmetrical_op_amp65 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_MainBias_1 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_2 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_3 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_4 outFirstStage outFirstStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_StageBias_6 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_Symmetrical_FirstStage_StageBias_7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Transconductor_8 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_Symmetrical_FirstStage_Transconductor_9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_StageBias_10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m_Symmetrical_SecondStage1_StageBias_11 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_Transconductor_12 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m_Symmetrical_SecondStage1_Transconductor_13 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_14 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_15 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_MainBias_17 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_18 ibias ibias sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_19 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_Symmetrical_SecondStage1_StageBias_20 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
.end symmetrical_op_amp65

