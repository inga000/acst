.suckt  two_stage_single_output_op_amp_125_1 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m3 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m4 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m5 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerOutputLoad2 sourcePmos sourcePmos pmos
m7 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerOutputLoad2 sourcePmos sourcePmos pmos
m9 sourceTransconductance outInputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c2 out sourceNmos 
m13 out outFirstStage sourceNmos sourceNmos nmos
m14 out ibias sourcePmos sourcePmos pmos
m15 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
m16 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m17 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m18 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_125_1

