** Name: two_stage_single_output_op_amp_10_9

.MACRO two_stage_single_output_op_amp_10_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=230e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=33e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=25e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=11e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=10e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=27e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=13e-6
mMainBias10 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=32e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=230e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=10e-6
mMainBias13 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=33e-6
mMainBias15 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=44e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=590e-6
mSimpleFirstStageLoad17 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=266e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.80001e-12
.EOM two_stage_single_output_op_amp_10_9

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 5.97901 mW
** Area: 10315 (mu_m)^2
** Transit frequency: 5.77001 MHz
** Transit frequency with error factor: 5.76358 MHz
** Slew rate: 9.12272 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** negPSRR: 105 dB
** posPSRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 1.76001 V
** VcmMax: 4.09001 V
** VcmMin: 0.960001 V


** Expected Currents: 
** NormalTransistorNmos: 1.38961e+07 muA
** NormalTransistorNmos: 6.34571e+07 muA
** NormalTransistorPmos: -5.64409e+07 muA
** DiodeTransistorPmos: -2.68039e+07 muA
** NormalTransistorPmos: -2.68039e+07 muA
** NormalTransistorPmos: -2.68039e+07 muA
** NormalTransistorNmos: 5.36051e+07 muA
** NormalTransistorNmos: 2.68031e+07 muA
** NormalTransistorNmos: 2.68031e+07 muA
** NormalTransistorNmos: 9.98418e+08 muA
** DiodeTransistorNmos: 9.98417e+08 muA
** NormalTransistorPmos: -9.98417e+08 muA
** DiodeTransistorNmos: 5.64401e+07 muA
** NormalTransistorNmos: 5.64391e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.38969e+07 muA
** DiodeTransistorPmos: -6.34579e+07 muA


** Expected Voltages: 
** ibias: 0.711001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.16201  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 1.08101  V
** outVoltageBiasXXpXX0: 3.73001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.40001  V
** out1: 3.83601  V
** sourceTransconductance: 1.84301  V
** inner: 1.07501  V


.END