** Name: one_stage_single_output_op_amp62

.MACRO one_stage_single_output_op_amp62 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=9e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=122e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=99e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=53e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=243e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=243e-6
mMainBias10 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad11 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=53e-6
mMainBias12 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=122e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=140e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=140e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=99e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageLoad18 out inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=8e-6 W=260e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp62

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 1.28101 mW
** Area: 6260 (mu_m)^2
** Transit frequency: 2.85701 MHz
** Transit frequency with error factor: 2.85692 MHz
** Slew rate: 3.82803 V/mu_s
** Phase margin: 88.2356°
** CMRR: 138 dB
** VoutMax: 4.45001 V
** VoutMin: 0.820001 V
** VcmMax: 3.06001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.76201e+06 muA
** NormalTransistorNmos: 1.00001e+07 muA
** NormalTransistorNmos: 7.68131e+07 muA
** NormalTransistorNmos: 1.15707e+08 muA
** NormalTransistorNmos: 7.68131e+07 muA
** NormalTransistorNmos: 1.15707e+08 muA
** DiodeTransistorPmos: -7.68139e+07 muA
** NormalTransistorPmos: -7.68139e+07 muA
** NormalTransistorPmos: -7.68139e+07 muA
** NormalTransistorPmos: -7.77889e+07 muA
** DiodeTransistorPmos: -7.77899e+07 muA
** NormalTransistorPmos: -3.88939e+07 muA
** NormalTransistorPmos: -3.88939e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -4.76299e+06 muA
** NormalTransistorPmos: -4.76399e+06 muA
** DiodeTransistorPmos: -1.00009e+07 muA


** Expected Voltages: 
** ibias: 1.18801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.68601  V
** out: 2.5  V
** outInputVoltageBiasXXpXX1: 3.27601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.13801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.61201  V
** out1: 4.24801  V
** sourceGCC1: 0.520001  V
** sourceGCC2: 0.520001  V
** sourceTransconductance: 3.27901  V
** inner: 4.13701  V


.END