** Name: two_stage_single_output_op_amp_46_7

.MACRO two_stage_single_output_op_amp_46_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=37e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=373e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=236e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=346e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=119e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=119e-6
mSecondStage1StageBias9 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=346e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=373e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=68e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=68e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=600e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=224e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=236e-6
mMainBias17 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=364e-6
mMainBias18 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=279e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.1001e-12
.EOM two_stage_single_output_op_amp_46_7

** Expected Performance Values: 
** Gain: 118 dB
** Power consumption: 8.94801 mW
** Area: 11286 (mu_m)^2
** Transit frequency: 3.96901 MHz
** Transit frequency with error factor: 3.96913 MHz
** Slew rate: 8.73727 V/mu_s
** Phase margin: 60.1606°
** CMRR: 139 dB
** VoutMax: 4.46001 V
** VoutMin: 0.150001 V
** VcmMax: 3.85001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -9.15589e+07 muA
** NormalTransistorPmos: -7.04729e+07 muA
** NormalTransistorNmos: 1.5061e+08 muA
** NormalTransistorNmos: 2.26652e+08 muA
** NormalTransistorNmos: 1.5061e+08 muA
** NormalTransistorNmos: 2.26652e+08 muA
** DiodeTransistorPmos: -1.50609e+08 muA
** DiodeTransistorPmos: -1.5061e+08 muA
** NormalTransistorPmos: -1.50609e+08 muA
** NormalTransistorPmos: -1.5061e+08 muA
** NormalTransistorPmos: -1.5208e+08 muA
** NormalTransistorPmos: -7.60409e+07 muA
** NormalTransistorPmos: -7.60409e+07 muA
** NormalTransistorNmos: 1.15432e+09 muA
** NormalTransistorPmos: -1.15431e+09 muA
** DiodeTransistorNmos: 9.15581e+07 muA
** DiodeTransistorNmos: 7.04721e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.89701  V
** outVoltageBiasXXnXX1: 0.915001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.28601  V
** innerTransistorStack2Load2: 4.28601  V
** out1: 3.53301  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.41601  V


.END