** Name: two_stage_single_output_op_amp_60_7

.MACRO two_stage_single_output_op_amp_60_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=189e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=82e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=77e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=33e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=33e-6
mSecondStage1StageBias9 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mFoldedCascodeFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=77e-6
mFoldedCascodeFirstStageLoad11 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=189e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=597e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=597e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=82e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=407e-6
mFoldedCascodeFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=233e-6
mMainBias18 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=142e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=31e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.5e-12
.EOM two_stage_single_output_op_amp_60_7

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 12.4601 mW
** Area: 14967 (mu_m)^2
** Transit frequency: 8.37801 MHz
** Transit frequency with error factor: 8.37787 MHz
** Slew rate: 7.6489 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.350001 V
** VcmMax: 3.03001 V
** VcmMin: -0.209999 V


** Expected Currents: 
** NormalTransistorPmos: -1.44684e+08 muA
** NormalTransistorPmos: -3.09609e+07 muA
** NormalTransistorNmos: 7.33291e+07 muA
** NormalTransistorNmos: 1.15105e+08 muA
** NormalTransistorNmos: 7.33291e+07 muA
** NormalTransistorNmos: 1.15105e+08 muA
** NormalTransistorPmos: -7.33299e+07 muA
** NormalTransistorPmos: -7.33299e+07 muA
** DiodeTransistorPmos: -7.33299e+07 muA
** NormalTransistorPmos: -8.35519e+07 muA
** DiodeTransistorPmos: -8.35509e+07 muA
** NormalTransistorPmos: -4.17759e+07 muA
** NormalTransistorPmos: -4.17759e+07 muA
** NormalTransistorNmos: 2.06622e+09 muA
** NormalTransistorPmos: -2.06621e+09 muA
** DiodeTransistorNmos: 1.44685e+08 muA
** DiodeTransistorNmos: 3.09601e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.19701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.10001  V
** outVoltageBiasXXnXX1: 1.10501  V
** outVoltageBiasXXnXX2: 0.755001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.07401  V
** out1: 3.32201  V
** sourceGCC1: 0.550001  V
** sourceGCC2: 0.550001  V
** sourceTransconductance: 3.22901  V
** inner: 4.09401  V


.END