.suckt  two_stage_fully_differential_op_amp_35_6 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 outInputVoltageBiasXXpXX3 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m4 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m5 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m6 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m7 outFeedback outFeedback sourceNmos sourceNmos nmos
m8 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m9 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m14 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m15 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m16 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m17 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m18 out1FirstStage ibias sourcePmos sourcePmos pmos
m19 out2FirstStage ibias sourcePmos sourcePmos pmos
m20 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m21 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m22 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m23 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m24 out1 outVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m25 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m26 out1 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m27 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m28 out2 outVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m29 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m30 out2 outInputVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos
m31 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m32 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m33 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m34 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m35 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m36 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m37 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m38 outInputVoltageBiasXXpXX3 outInputVoltageBiasXXpXX3 VoltageBiasXXpXX3Yinner VoltageBiasXXpXX3Yinner pmos
m39 VoltageBiasXXpXX3Yinner outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m40 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_35_6

