** Name: symmetrical_op_amp50

.MACRO symmetrical_op_amp50 ibias in1 in2 out sourceNmos sourcePmos
m1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=20e-6
m2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=37e-6
m3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=37e-6
m4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=19e-6
m5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=98e-6
m6 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=2e-6 W=10e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=44e-6
m8 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=3e-6 W=5e-6
m9 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=5e-6
m10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=110e-6
m11 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=110e-6
m12 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=448e-6
m13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=53e-6
m14 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=8e-6
m15 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=53e-6
m16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=44e-6
m17 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=98e-6
m18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp50

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 1.75701 mW
** Area: 4216 (mu_m)^2
** Transit frequency: 3.53001 MHz
** Transit frequency with error factor: 3.52992 MHz
** Slew rate: 3.50001 V/mu_s
** Phase margin: 61.3065°
** CMRR: 142 dB
** negPSRR: 44 dB
** posPSRR: 46 dB
** VoutMax: 3.54001 V
** VoutMin: 0.650001 V
** VcmMax: 3.12001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorPmos: -2.37884e+08 muA
** DiodeTransistorNmos: 1.17551e+07 muA
** DiodeTransistorNmos: 1.17551e+07 muA
** NormalTransistorPmos: -2.35109e+07 muA
** DiodeTransistorPmos: -2.35099e+07 muA
** NormalTransistorPmos: -1.17559e+07 muA
** NormalTransistorPmos: -1.17559e+07 muA
** NormalTransistorNmos: 3.50041e+07 muA
** NormalTransistorNmos: 3.50031e+07 muA
** NormalTransistorPmos: -3.50049e+07 muA
** NormalTransistorPmos: -3.50059e+07 muA
** DiodeTransistorPmos: -3.49209e+07 muA
** DiodeTransistorPmos: -3.49219e+07 muA
** NormalTransistorNmos: 3.49201e+07 muA
** NormalTransistorNmos: 3.49191e+07 muA
** DiodeTransistorNmos: 2.37885e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.27301  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 1.05101  V
** inSourceStageBiasComplementarySecondStage: 4.23601  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 3.04401  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.13801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.22101  V
** innerStageBias: 4.30501  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V
** inner: 4.13301  V


.END