** Name: two_stage_single_output_op_amp_12_10

.MACRO two_stage_single_output_op_amp_12_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias2 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mSimpleFirstStageTransconductor3 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=140e-6
mSimpleFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=43e-6
mSecondStage1StageBias5 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=472e-6
mSimpleFirstStageTransconductor6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=140e-6
mMainBias7 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=162e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=49e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=49e-6
mSimpleFirstStageLoad10 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=103e-6
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=373e-6
mSecondStage1Transconductor12 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad13 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=103e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.2001e-12
.EOM two_stage_single_output_op_amp_12_10

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 8.51101 mW
** Area: 5054 (mu_m)^2
** Transit frequency: 6.55501 MHz
** Transit frequency with error factor: 6.55179 MHz
** Slew rate: 6.17795 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 109 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 0.300001 V
** VcmMax: 4.91001 V
** VcmMin: 0.850001 V


** Expected Currents: 
** NormalTransistorNmos: 4.06136e+08 muA
** NormalTransistorPmos: -5.33309e+07 muA
** NormalTransistorPmos: -5.33319e+07 muA
** NormalTransistorPmos: -5.33309e+07 muA
** NormalTransistorPmos: -5.33319e+07 muA
** NormalTransistorNmos: 1.0666e+08 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 1.17942e+09 muA
** NormalTransistorPmos: -1.17941e+09 muA
** NormalTransistorPmos: -1.17941e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.06135e+08 muA


** Expected Voltages: 
** ibias: 0.702001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.01601  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.42001  V
** innerTransistorStack2Load1: 4.42001  V
** out1: 3.94001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.58001  V


.END