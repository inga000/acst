.suckt  two_stage_fully_differential_op_amp_44_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m4 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m5 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m6 outFeedback outFeedback sourceNmos sourceNmos nmos
m7 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m8 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m9 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m10 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m11 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m15 out1FirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m16 out2FirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m17 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m18 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m19 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m20 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m21 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m22 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m23 out1 outVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m24 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m25 out1 ibias SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m26 SecondStage1YinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m27 out2 outVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m28 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m29 out2 ibias SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m30 SecondStage2YinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m31 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m32 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m33 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m34 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m35 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos
m36 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos
m37 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_44_4

