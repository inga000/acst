** Name: symmetrical_op_amp196

.MACRO symmetrical_op_amp196 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=10e-6
mSecondStage1StageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=16e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=2e-6 W=16e-6
mSymmetricalFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=92e-6
mMainBias5 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=92e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias7 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=16e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=10e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=93e-6
mSecondStage1StageBias10 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=2e-6 W=16e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=93e-6
mMainBias12 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=100e-6
mSymmetricalFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=49e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=49e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=72e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=72e-6
mSymmetricalFirstStageLoad17 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=112e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=166e-6
mSecondStage1Transconductor19 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=166e-6
mSymmetricalFirstStageLoad20 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=112e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp196

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 1.67101 mW
** Area: 4652 (mu_m)^2
** Transit frequency: 6.95801 MHz
** Transit frequency with error factor: 6.95806 MHz
** Slew rate: 6.67072 V/mu_s
** Phase margin: 73.3387°
** CMRR: 141 dB
** negPSRR: 130 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 1.03001 V
** VcmMax: 4.81001 V
** VcmMin: 1.44001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00151e+08 muA
** NormalTransistorPmos: -4.51569e+07 muA
** NormalTransistorPmos: -4.51579e+07 muA
** NormalTransistorPmos: -4.51569e+07 muA
** NormalTransistorPmos: -4.51579e+07 muA
** NormalTransistorNmos: 9.03131e+07 muA
** DiodeTransistorNmos: 9.03141e+07 muA
** NormalTransistorNmos: 4.51561e+07 muA
** NormalTransistorNmos: 4.51561e+07 muA
** NormalTransistorNmos: 6.68381e+07 muA
** DiodeTransistorNmos: 6.68371e+07 muA
** NormalTransistorPmos: -6.68389e+07 muA
** NormalTransistorPmos: -6.68379e+07 muA
** DiodeTransistorNmos: 6.68381e+07 muA
** NormalTransistorNmos: 6.68371e+07 muA
** NormalTransistorPmos: -6.68389e+07 muA
** NormalTransistorPmos: -6.68379e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.0015e+08 muA


** Expected Voltages: 
** ibias: 1.29201  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 0.718001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 1.43601  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.647001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94301  V
** innerTransconductance: 4.40001  V
** inner: 0.716001  V
** inner: 4.40001  V
** inner: 0.643001  V


.END