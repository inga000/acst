** Name: two_stage_single_output_op_amp_189_9

.MACRO two_stage_single_output_op_amp_189_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=9e-6 W=9e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=13e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=168e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=30e-6
m5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=23e-6
m6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=112e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=13e-6
m8 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=168e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=10e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=10e-6
m11 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=77e-6
m12 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=23e-6
m13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=10e-6
m14 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=9e-6 W=12e-6
m15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
m16 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=204e-6
m17 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=9e-6
m18 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=596e-6
m19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=67e-6
m20 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=112e-6
m21 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=112e-6
m22 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=7e-6 W=596e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_189_9

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 4.72601 mW
** Area: 14611 (mu_m)^2
** Transit frequency: 3.38801 MHz
** Transit frequency with error factor: 3.38587 MHz
** Slew rate: 3.77233 V/mu_s
** Phase margin: 65.3172°
** CMRR: 112 dB
** VoutMax: 4.25 V
** VoutMin: 1.16001 V
** VcmMax: 4.62001 V
** VcmMin: 1.54001 V


** Expected Currents: 
** NormalTransistorPmos: -5.24439e+07 muA
** NormalTransistorPmos: -6.90699e+06 muA
** NormalTransistorNmos: 7.88221e+07 muA
** NormalTransistorNmos: 7.88211e+07 muA
** DiodeTransistorNmos: 7.88221e+07 muA
** NormalTransistorPmos: -8.76829e+07 muA
** NormalTransistorPmos: -8.76819e+07 muA
** NormalTransistorPmos: -8.76829e+07 muA
** NormalTransistorPmos: -8.76819e+07 muA
** NormalTransistorNmos: 1.77211e+07 muA
** NormalTransistorNmos: 1.77201e+07 muA
** NormalTransistorNmos: 8.86101e+06 muA
** NormalTransistorNmos: 8.86101e+06 muA
** NormalTransistorNmos: 6.90431e+08 muA
** DiodeTransistorNmos: 6.9043e+08 muA
** NormalTransistorPmos: -6.9043e+08 muA
** DiodeTransistorNmos: 5.24431e+07 muA
** NormalTransistorNmos: 5.24441e+07 muA
** DiodeTransistorNmos: 6.90601e+06 muA
** DiodeTransistorNmos: 6.90501e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.25101  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.57001  V
** outSourceVoltageBiasXXnXX1: 0.785001  V
** outSourceVoltageBiasXXnXX2: 0.561001  V
** outSourceVoltageBiasXXpXX1: 3.88501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.940001  V
** innerStageBias: 0.448001  V
** innerTransistorStack1Load2: 3.93701  V
** innerTransistorStack2Load2: 3.93701  V
** out1: 2.09501  V
** sourceTransconductance: 1.91701  V
** inner: 0.786001  V


.END