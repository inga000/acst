** Name: two_stage_single_output_op_amp_45_7

.MACRO two_stage_single_output_op_amp_45_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=163e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=186e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=42e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=52e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=83e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=286e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=286e-6
mMainBias9 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=116e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=529e-6
mFoldedCascodeFirstStageLoad11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=83e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=186e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=86e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=86e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=554e-6
mMainBias16 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=153e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=494e-6
mFoldedCascodeFirstStageLoad18 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=421e-6
mMainBias19 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=437e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.30001e-12
.EOM two_stage_single_output_op_amp_45_7

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 4.66701 mW
** Area: 14259 (mu_m)^2
** Transit frequency: 5.39401 MHz
** Transit frequency with error factor: 5.39382 MHz
** Slew rate: 11.3806 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 4.80001 V
** VoutMin: 0.150001 V
** VcmMax: 3.79001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 7.43891e+07 muA
** NormalTransistorPmos: -3.64359e+07 muA
** NormalTransistorPmos: -1.03485e+08 muA
** NormalTransistorNmos: 1.14875e+08 muA
** NormalTransistorNmos: 1.81576e+08 muA
** NormalTransistorNmos: 1.14874e+08 muA
** NormalTransistorNmos: 1.81576e+08 muA
** DiodeTransistorPmos: -1.14875e+08 muA
** NormalTransistorPmos: -1.14873e+08 muA
** NormalTransistorPmos: -1.14875e+08 muA
** NormalTransistorPmos: -1.33401e+08 muA
** NormalTransistorPmos: -6.67009e+07 muA
** NormalTransistorPmos: -6.67009e+07 muA
** NormalTransistorNmos: 3.3585e+08 muA
** NormalTransistorPmos: -3.35849e+08 muA
** DiodeTransistorNmos: 3.64351e+07 muA
** DiodeTransistorNmos: 1.03486e+08 muA
** DiodeTransistorPmos: -7.43899e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.20501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.976001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.24001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.57601  V
** out1: 4.25  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.47901  V


.END