** Name: two_stage_single_output_op_amp_54_1

.MACRO two_stage_single_output_op_amp_54_1 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
m2 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=11e-6
m3 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=89e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=25e-6
m5 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=211e-6
m6 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=55e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=491e-6
m8 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=140e-6
m9 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=55e-6
m10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=352e-6
m11 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=352e-6
m12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=79e-6
m13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=79e-6
m14 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=9e-6 W=164e-6
m15 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=136e-6
m16 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=551e-6
m17 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=590e-6
m18 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=551e-6
m19 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=89e-6
m20 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=89e-6
Capacitor1 outFirstStage out 21e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_54_1

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 11.1641 mW
** Area: 14275 (mu_m)^2
** Transit frequency: 6.09701 MHz
** Transit frequency with error factor: 6.09731 MHz
** Slew rate: 5.29925 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.66001 V
** VoutMin: 0.300001 V
** VcmMax: 5.06001 V
** VcmMin: 0.900001 V


** Expected Currents: 
** NormalTransistorNmos: 1.26917e+08 muA
** NormalTransistorNmos: 1.89002e+08 muA
** NormalTransistorPmos: -2.83477e+08 muA
** NormalTransistorPmos: -1.11889e+08 muA
** NormalTransistorPmos: -1.85274e+08 muA
** NormalTransistorPmos: -1.11889e+08 muA
** NormalTransistorPmos: -1.85274e+08 muA
** NormalTransistorNmos: 1.1189e+08 muA
** NormalTransistorNmos: 1.11889e+08 muA
** NormalTransistorNmos: 1.1189e+08 muA
** NormalTransistorNmos: 1.11889e+08 muA
** NormalTransistorNmos: 1.46769e+08 muA
** NormalTransistorNmos: 7.33841e+07 muA
** NormalTransistorNmos: 7.33841e+07 muA
** NormalTransistorNmos: 1.25294e+09 muA
** NormalTransistorPmos: -1.25293e+09 muA
** DiodeTransistorNmos: 2.83478e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.26916e+08 muA
** DiodeTransistorPmos: -1.89001e+08 muA


** Expected Voltages: 
** ibias: 0.715001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.910001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outVoltageBiasXXpXX2: 4.09301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.350001  V
** innerTransistorStack2Load2: 0.350001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.91301  V


.END