** Name: two_stage_single_output_op_amp_59_7

.MACRO two_stage_single_output_op_amp_59_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=94e-6
m3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=592e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
m7 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=371e-6
m8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=371e-6
m9 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=137e-6
m10 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=137e-6
m11 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=411e-6
m12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=600e-6
m13 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
m14 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=283e-6
m15 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=337e-6
m16 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=592e-6
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=404e-6
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=404e-6
m19 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=574e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 14.4001e-12
.EOM two_stage_single_output_op_amp_59_7

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 14.9781 mW
** Area: 13931 (mu_m)^2
** Transit frequency: 7.96701 MHz
** Transit frequency with error factor: 7.96643 MHz
** Slew rate: 16.5394 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 4.5 V
** VoutMin: 0.190001 V
** VcmMax: 3 V
** VcmMin: -0.369999 V


** Expected Currents: 
** NormalTransistorPmos: -4.15689e+07 muA
** NormalTransistorPmos: -2.81422e+08 muA
** NormalTransistorNmos: 2.42414e+08 muA
** NormalTransistorNmos: 4.10158e+08 muA
** NormalTransistorNmos: 2.42414e+08 muA
** NormalTransistorNmos: 4.10158e+08 muA
** NormalTransistorPmos: -2.42413e+08 muA
** NormalTransistorPmos: -2.42413e+08 muA
** DiodeTransistorPmos: -2.42413e+08 muA
** NormalTransistorPmos: -3.3549e+08 muA
** NormalTransistorPmos: -3.35491e+08 muA
** NormalTransistorPmos: -1.67744e+08 muA
** NormalTransistorPmos: -1.67744e+08 muA
** NormalTransistorNmos: 1.83235e+09 muA
** NormalTransistorPmos: -1.83234e+09 muA
** DiodeTransistorNmos: 4.15681e+07 muA
** DiodeTransistorNmos: 2.81423e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.93501  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.946001  V
** outVoltageBiasXXnXX2: 0.594001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.28501  V
** innerStageBias: 4.14201  V
** out1: 3.57101  V
** sourceGCC1: 0.389001  V
** sourceGCC2: 0.389001  V
** sourceTransconductance: 3.51901  V


.END