** Name: two_stage_single_output_op_amp_205_12

.MACRO two_stage_single_output_op_amp_205_12 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=5e-6 W=39e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=39e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=8e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=4e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=425e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=38e-6
mSimpleFirstStageTransconductor9 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=124e-6
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=248e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=9e-6 W=39e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=73e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=425e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=39e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=124e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=574e-6
mMainBias18 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=39e-6
mSimpleFirstStageLoad19 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=389e-6
mSimpleFirstStageLoad20 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=533e-6
mSimpleFirstStageLoad21 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=533e-6
mSecondStage1Transconductor22 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=552e-6
mSecondStage1Transconductor23 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad24 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=389e-6
mMainBias25 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=28e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.7001e-12
.EOM two_stage_single_output_op_amp_205_12

** Expected Performance Values: 
** Gain: 141 dB
** Power consumption: 11.4321 mW
** Area: 14995 (mu_m)^2
** Transit frequency: 6.00701 MHz
** Transit frequency with error factor: 6.00519 MHz
** Slew rate: 5.6619 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** VoutMax: 4.25 V
** VoutMin: 1.10001 V
** VcmMax: 4.88001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorNmos: 2.74142e+08 muA
** NormalTransistorNmos: 1.87571e+07 muA
** NormalTransistorPmos: -1.37289e+07 muA
** DiodeTransistorNmos: 2.00496e+08 muA
** NormalTransistorNmos: 2.00497e+08 muA
** NormalTransistorNmos: 2.00496e+08 muA
** DiodeTransistorNmos: 2.00497e+08 muA
** NormalTransistorPmos: -2.59539e+08 muA
** NormalTransistorPmos: -2.5954e+08 muA
** NormalTransistorPmos: -2.59539e+08 muA
** NormalTransistorPmos: -2.5954e+08 muA
** NormalTransistorNmos: 1.18088e+08 muA
** NormalTransistorNmos: 1.18088e+08 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorNmos: 1.45079e+09 muA
** DiodeTransistorNmos: 1.45079e+09 muA
** NormalTransistorPmos: -1.45078e+09 muA
** NormalTransistorPmos: -1.45078e+09 muA
** DiodeTransistorNmos: 1.37281e+07 muA
** NormalTransistorNmos: 1.37271e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.74141e+08 muA
** DiodeTransistorPmos: -1.87579e+07 muA


** Expected Voltages: 
** ibias: 1.20201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.05201  V
** outInputVoltageBiasXXnXX1: 1.50401  V
** outSourceVoltageBiasXXnXX1: 0.752001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.10501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.10601  V
** innerStageBias: 0.520001  V
** innerTransistorStack1Load1: 1.14801  V
** innerTransistorStack1Load2: 4.44301  V
** innerTransistorStack2Load1: 1.14801  V
** innerTransistorStack2Load2: 4.44301  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.61601  V
** inner: 0.749001  V


.END