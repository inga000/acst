** Name: two_stage_single_output_op_amp_62_9

.MACRO two_stage_single_output_op_amp_62_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=8e-6 W=140e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=17e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=296e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=68e-6
m5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=89e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=300e-6
m7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=6e-6
m8 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=48e-6
m9 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=296e-6
m10 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=8e-6 W=71e-6
m11 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=33e-6
m12 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=8e-6 W=71e-6
m13 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=68e-6
m14 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=68e-6
m15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=17e-6
m16 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=359e-6
m17 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=390e-6
m18 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=134e-6
m19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=287e-6
m20 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=48e-6
m21 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=15e-6
m22 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=15e-6
m23 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=300e-6
m24 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=89e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_62_9

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 3.79701 mW
** Area: 14900 (mu_m)^2
** Transit frequency: 2.73601 MHz
** Transit frequency with error factor: 2.73647 MHz
** Slew rate: 5.2743 V/mu_s
** Phase margin: 68.755°
** CMRR: 131 dB
** VoutMax: 4.60001 V
** VoutMin: 0.700001 V
** VcmMax: 3.04001 V
** VcmMin: -0.319999 V


** Expected Currents: 
** NormalTransistorNmos: 2.01471e+07 muA
** NormalTransistorPmos: -3.23799e+07 muA
** NormalTransistorPmos: -4.06939e+07 muA
** NormalTransistorNmos: 2.40231e+07 muA
** NormalTransistorNmos: 4.11841e+07 muA
** NormalTransistorNmos: 2.40201e+07 muA
** NormalTransistorNmos: 4.11791e+07 muA
** DiodeTransistorPmos: -2.40219e+07 muA
** NormalTransistorPmos: -2.40209e+07 muA
** NormalTransistorPmos: -2.40219e+07 muA
** NormalTransistorPmos: -3.43189e+07 muA
** DiodeTransistorPmos: -3.43179e+07 muA
** NormalTransistorPmos: -1.71599e+07 muA
** NormalTransistorPmos: -1.71599e+07 muA
** NormalTransistorNmos: 5.63771e+08 muA
** DiodeTransistorNmos: 5.63771e+08 muA
** NormalTransistorPmos: -5.6377e+08 muA
** DiodeTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** DiodeTransistorNmos: 4.06931e+07 muA
** DiodeTransistorNmos: 4.06941e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -2.01479e+07 muA


** Expected Voltages: 
** ibias: 3.48101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.21401  V
** out: 2.5  V
** outFirstStage: 4.03201  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.644001  V
** outSourceVoltageBiasXXpXX1: 4.24101  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.42301  V
** out1: 4.14501  V
** sourceGCC1: 0.630001  V
** sourceGCC2: 0.630001  V
** sourceTransconductance: 3.50101  V
** inner: 0.555001  V
** inner: 4.23901  V


.END