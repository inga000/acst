** Name: two_stage_single_output_op_amp_34_12

.MACRO two_stage_single_output_op_amp_34_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=8e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=256e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=110e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=372e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=61e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=37e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=52e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=61e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=110e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=256e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mSecondStage1StageBias12 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=372e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=61e-6
mMainBias14 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=142e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=61e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=578e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=308e-6
mSimpleFirstStageLoad19 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=13e-6
mMainBias20 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=86e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_34_12

** Expected Performance Values: 
** Gain: 145 dB
** Power consumption: 3.77001 mW
** Area: 14910 (mu_m)^2
** Transit frequency: 6.06401 MHz
** Transit frequency with error factor: 6.06146 MHz
** Slew rate: 5.715 V/mu_s
** Phase margin: 64.1713°
** CMRR: 103 dB
** negPSRR: 109 dB
** posPSRR: 98 dB
** VoutMax: 4.29001 V
** VoutMin: 0.890001 V
** VcmMax: 4.09001 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorNmos: 2.60941e+07 muA
** NormalTransistorNmos: 1.75992e+08 muA
** NormalTransistorPmos: -5.95149e+07 muA
** DiodeTransistorPmos: -1.29109e+07 muA
** NormalTransistorPmos: -1.29109e+07 muA
** NormalTransistorPmos: -1.29109e+07 muA
** NormalTransistorNmos: 2.58191e+07 muA
** DiodeTransistorNmos: 2.58181e+07 muA
** NormalTransistorNmos: 1.29101e+07 muA
** NormalTransistorNmos: 1.29101e+07 muA
** NormalTransistorNmos: 4.56478e+08 muA
** DiodeTransistorNmos: 4.56479e+08 muA
** NormalTransistorPmos: -4.56477e+08 muA
** NormalTransistorPmos: -4.56478e+08 muA
** DiodeTransistorNmos: 5.95141e+07 muA
** NormalTransistorNmos: 5.95141e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.60949e+07 muA
** DiodeTransistorPmos: -1.75991e+08 muA


** Expected Voltages: 
** ibias: 1.29201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.22501  V
** outInputVoltageBiasXXnXX1: 1.12601  V
** outSourceVoltageBiasXXnXX1: 0.563001  V
** outSourceVoltageBiasXXnXX2: 0.647001  V
** outVoltageBiasXXpXX0: 3.99401  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.65701  V
** out1: 4.09301  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.74701  V
** inner: 0.563001  V
** inner: 0.643001  V


.END