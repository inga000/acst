** Name: one_stage_single_output_op_amp124

.MACRO one_stage_single_output_op_amp124 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=19e-6
mTelescopicFirstStageStageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=238e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=37e-6
mTelescopicFirstStageLoad4 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=40e-6
mTelescopicFirstStageLoad5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=10e-6
mTelescopicFirstStageLoad7 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=56e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=28e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=2e-6 W=28e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=19e-6
mMainBias11 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=19e-6
mTelescopicFirstStageLoad12 out outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=56e-6
mTelescopicFirstStageStageBias13 sourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=238e-6
mTelescopicFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=40e-6
mTelescopicFirstStageLoad15 out FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=40e-6
mMainBias16 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=70e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp124

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 0.718001 mW
** Area: 4333 (mu_m)^2
** Transit frequency: 2.82501 MHz
** Transit frequency with error factor: 2.82486 MHz
** Slew rate: 6.1693 V/mu_s
** Phase margin: 87.0896°
** CMRR: 146 dB
** VoutMax: 4.05001 V
** VoutMin: 1.06001 V
** VcmMax: 3.74001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00641e+07 muA
** NormalTransistorPmos: -7.02469e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** DiodeTransistorPmos: -2.66659e+07 muA
** NormalTransistorPmos: -2.66669e+07 muA
** NormalTransistorPmos: -2.66659e+07 muA
** DiodeTransistorPmos: -2.66669e+07 muA
** NormalTransistorNmos: 1.23578e+08 muA
** DiodeTransistorNmos: 1.23579e+08 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 7.02461e+07 muA
** DiodeTransistorPmos: -1.00649e+07 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.68301  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.581001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerOutputLoad2: 3.48401  V
** innerSourceLoad2: 4.24201  V
** innerTransistorStack1Load2: 4.24101  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.579001  V


.END