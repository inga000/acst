** Name: symmetrical_op_amp36

.MACRO symmetrical_op_amp36 ibias in1 in2 out sourceNmos sourcePmos
m1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
m2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=133e-6
m3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=133e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
m5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=395e-6
m6 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=6e-6 W=147e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m8 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=3e-6 W=93e-6
m9 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=93e-6
m10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=129e-6
m11 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=129e-6
m12 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=35e-6
m13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=403e-6
m14 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=6e-6 W=182e-6
m15 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=403e-6
m16 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=503e-6
m17 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=252e-6
m18 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=395e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp36

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 5.29701 mW
** Area: 9430 (mu_m)^2
** Transit frequency: 20.8531 MHz
** Transit frequency with error factor: 20.8528 MHz
** Slew rate: 24.4924 V/mu_s
** Phase margin: 80.7871°
** CMRR: 142 dB
** negPSRR: 47 dB
** posPSRR: 51 dB
** VoutMax: 3.31001 V
** VoutMin: 0.460001 V
** VcmMax: 3.11001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorPmos: -3.54849e+07 muA
** DiodeTransistorNmos: 2.54991e+08 muA
** DiodeTransistorNmos: 2.54991e+08 muA
** NormalTransistorPmos: -5.0998e+08 muA
** NormalTransistorPmos: -5.09979e+08 muA
** NormalTransistorPmos: -2.5499e+08 muA
** NormalTransistorPmos: -2.5499e+08 muA
** NormalTransistorNmos: 2.45699e+08 muA
** NormalTransistorNmos: 2.45698e+08 muA
** NormalTransistorPmos: -2.45698e+08 muA
** NormalTransistorPmos: -2.45699e+08 muA
** DiodeTransistorPmos: -2.48179e+08 muA
** DiodeTransistorPmos: -2.4818e+08 muA
** NormalTransistorNmos: 2.4818e+08 muA
** NormalTransistorNmos: 2.48179e+08 muA
** DiodeTransistorNmos: 3.54841e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.861001  V
** inSourceStageBiasComplementarySecondStage: 3.97701  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 2.66301  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.29701  V
** sourceTransconductance: 3.25201  V
** innerStageBias: 3.89701  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END