.suckt  two_stage_fully_differential_op_amp_2_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_3 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_Load_5 outFeedback outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_6 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_8 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackStage_Transconductor_10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FeedbackStage_Transconductor_13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FirstStage_Load_14 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_15 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_StageBias_16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Transconductor_17 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_FullyDifferential_FirstStage_Transconductor_18 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_Transconductor_19 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m_FullyDifferential_SecondStage1_Transconductor_20 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_21 out1 outVoltageBiasXXpXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m_FullyDifferential_SecondStage1_StageBias_22 SecondStage1YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_Transconductor_23 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m_FullyDifferential_SecondStage2_Transconductor_24 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_StageBias_25 out2 outVoltageBiasXXpXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m_FullyDifferential_SecondStage2_StageBias_26 SecondStage2YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_27 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_28 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_29 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_30 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_2_4

