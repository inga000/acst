** Name: two_stage_single_output_op_amp_37_8

.MACRO two_stage_single_output_op_amp_37_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=8e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mSimpleFirstStageStageBias4 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=89e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=62e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=29e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mMainBias8 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=46e-6
mSecondStage1StageBias9 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=178e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=62e-6
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=76e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=76e-6
mSimpleFirstStageLoad13 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=123e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=542e-6
mSimpleFirstStageLoad15 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=123e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_37_8

** Expected Performance Values: 
** Gain: 105 dB
** Power consumption: 2.49901 mW
** Area: 4741 (mu_m)^2
** Transit frequency: 6.84301 MHz
** Transit frequency with error factor: 6.839 MHz
** Slew rate: 6.44925 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** negPSRR: 121 dB
** posPSRR: 105 dB
** VoutMax: 4.80001 V
** VoutMin: 0.840001 V
** VcmMax: 5.20001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 3.04591e+07 muA
** NormalTransistorPmos: -2.95229e+07 muA
** NormalTransistorPmos: -2.95239e+07 muA
** NormalTransistorPmos: -2.95229e+07 muA
** NormalTransistorPmos: -2.95239e+07 muA
** NormalTransistorNmos: 5.90431e+07 muA
** NormalTransistorNmos: 5.90421e+07 muA
** NormalTransistorNmos: 2.95221e+07 muA
** NormalTransistorNmos: 2.95221e+07 muA
** NormalTransistorNmos: 4.00319e+08 muA
** NormalTransistorNmos: 4.00318e+08 muA
** NormalTransistorPmos: -4.00318e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.04599e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.23201  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.499001  V
** innerTransistorStack1Load1: 4.41401  V
** innerTransistorStack2Load1: 4.41401  V
** out1: 4.22701  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.485001  V


.END