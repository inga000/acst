** Name: two_stage_single_output_op_amp_76_9

.MACRO two_stage_single_output_op_amp_76_9 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=103e-6
m2 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=5e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=31e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=362e-6
m5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=6e-6 W=29e-6
m6 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=22e-6
m7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=42e-6
m8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=22e-6
m9 outFirstStage outVoltageBiasXXnXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=26e-6
m10 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=362e-6
m11 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=22e-6
m12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=5e-6
m13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=5e-6
m14 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=31e-6
m15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=103e-6
m16 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=56e-6
m18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=205e-6
m19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=129e-6
m20 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=62e-6
m21 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=395e-6
m22 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=56e-6
m23 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=54e-6
m24 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=54e-6
Capacitor1 outFirstStage out 4.5e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_76_9

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 12.1051 mW
** Area: 7731 (mu_m)^2
** Transit frequency: 3.07801 MHz
** Transit frequency with error factor: 3.07752 MHz
** Slew rate: 3.52063 V/mu_s
** Phase margin: 74.4846°
** CMRR: 137 dB
** VoutMax: 4.25 V
** VoutMin: 1.14001 V
** VcmMax: 5.09001 V
** VcmMin: 1.45001 V


** Expected Currents: 
** NormalTransistorPmos: -5.96089e+07 muA
** NormalTransistorPmos: -2.86489e+07 muA
** NormalTransistorPmos: -1.81303e+08 muA
** NormalTransistorPmos: -1.59199e+07 muA
** NormalTransistorPmos: -2.49529e+07 muA
** NormalTransistorPmos: -1.59199e+07 muA
** NormalTransistorPmos: -2.49529e+07 muA
** DiodeTransistorNmos: 1.59191e+07 muA
** NormalTransistorNmos: 1.59191e+07 muA
** NormalTransistorNmos: 1.59191e+07 muA
** NormalTransistorNmos: 1.80631e+07 muA
** DiodeTransistorNmos: 1.80621e+07 muA
** NormalTransistorNmos: 9.03201e+06 muA
** NormalTransistorNmos: 9.03201e+06 muA
** NormalTransistorNmos: 2.08145e+09 muA
** DiodeTransistorNmos: 2.08145e+09 muA
** NormalTransistorPmos: -2.08144e+09 muA
** DiodeTransistorNmos: 5.96081e+07 muA
** NormalTransistorNmos: 5.96071e+07 muA
** DiodeTransistorNmos: 2.86481e+07 muA
** NormalTransistorNmos: 2.86471e+07 muA
** DiodeTransistorNmos: 1.81304e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.24801  V
** outInputVoltageBiasXXnXX2: 1.54401  V
** outSourceVoltageBiasXXnXX1: 0.624001  V
** outSourceVoltageBiasXXnXX2: 0.772001  V
** outSourceVoltageBiasXXpXX1: 4.11601  V
** outVoltageBiasXXnXX3: 1.07401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.461001  V
** out1: 0.666001  V
** sourceGCC1: 4.13701  V
** sourceGCC2: 4.13701  V
** sourceTransconductance: 1.88801  V
** inner: 0.624001  V
** inner: 0.770001  V


.END