** Name: two_stage_single_output_op_amp_188_8

.MACRO two_stage_single_output_op_amp_188_8 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=24e-6
m2 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=31e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=53e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=17e-6
m5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
m6 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=31e-6
m7 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=319e-6
m8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=4e-6
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=48e-6
m10 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
m11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=48e-6
m12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=53e-6
m13 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=271e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=24e-6
m15 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=469e-6
m16 outFirstStage ibias sourcePmos sourcePmos pmos4 L=4e-6 W=161e-6
m17 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=51e-6
m18 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=180e-6
m19 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=161e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.70001e-12
.EOM two_stage_single_output_op_amp_188_8

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 5.77001 mW
** Area: 7299 (mu_m)^2
** Transit frequency: 3.97901 MHz
** Transit frequency with error factor: 3.96959 MHz
** Slew rate: 3.75019 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 0.800001 V
** VcmMax: 5.14001 V
** VcmMin: 1.5 V


** Expected Currents: 
** NormalTransistorPmos: -1.66239e+07 muA
** NormalTransistorPmos: -5.90449e+07 muA
** NormalTransistorNmos: 3.46521e+07 muA
** NormalTransistorNmos: 3.46511e+07 muA
** DiodeTransistorNmos: 3.46521e+07 muA
** NormalTransistorPmos: -5.29369e+07 muA
** NormalTransistorPmos: -5.29369e+07 muA
** NormalTransistorNmos: 3.65691e+07 muA
** DiodeTransistorNmos: 3.65681e+07 muA
** NormalTransistorNmos: 1.82851e+07 muA
** NormalTransistorNmos: 1.82851e+07 muA
** NormalTransistorNmos: 9.52389e+08 muA
** NormalTransistorNmos: 9.52388e+08 muA
** NormalTransistorPmos: -9.52388e+08 muA
** DiodeTransistorNmos: 1.66231e+07 muA
** NormalTransistorNmos: 1.66221e+07 muA
** DiodeTransistorNmos: 5.90441e+07 muA
** DiodeTransistorNmos: 5.90431e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.16601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.35001  V
** outInputVoltageBiasXXnXX2: 1.16301  V
** outSourceVoltageBiasXXnXX1: 0.675001  V
** outSourceVoltageBiasXXnXX2: 0.608001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.04801  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.570001  V
** inner: 0.673001  V


.END