** Name: two_stage_single_output_op_amp_65_8

.MACRO two_stage_single_output_op_amp_65_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=11e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=40e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=224e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=224e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=600e-6
mMainBias9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=158e-6
mMainBias10 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=70e-6
mSecondStage1StageBias11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=6e-6 W=456e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=40e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=113e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=87e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=87e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=109e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=30e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=30e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=99e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=372e-6
mFoldedCascodeFirstStageLoad21 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=109e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.8001e-12
.EOM two_stage_single_output_op_amp_65_8

** Expected Performance Values: 
** Gain: 134 dB
** Power consumption: 2.10801 mW
** Area: 12222 (mu_m)^2
** Transit frequency: 2.81301 MHz
** Transit frequency with error factor: 2.81339 MHz
** Slew rate: 3.6847 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 4.83001 V
** VoutMin: 0.730001 V
** VcmMax: 3.34001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 5.13391e+07 muA
** NormalTransistorNmos: 2.25491e+07 muA
** NormalTransistorNmos: 4.73161e+07 muA
** NormalTransistorNmos: 7.13441e+07 muA
** NormalTransistorNmos: 4.73161e+07 muA
** NormalTransistorNmos: 7.13441e+07 muA
** NormalTransistorPmos: -4.73169e+07 muA
** NormalTransistorPmos: -4.73179e+07 muA
** NormalTransistorPmos: -4.73169e+07 muA
** NormalTransistorPmos: -4.73179e+07 muA
** NormalTransistorPmos: -4.80589e+07 muA
** NormalTransistorPmos: -4.80599e+07 muA
** NormalTransistorPmos: -2.40289e+07 muA
** NormalTransistorPmos: -2.40289e+07 muA
** NormalTransistorNmos: 1.94962e+08 muA
** NormalTransistorNmos: 1.94961e+08 muA
** NormalTransistorPmos: -1.94961e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.13399e+07 muA
** DiodeTransistorPmos: -2.25499e+07 muA


** Expected Voltages: 
** ibias: 1.21401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.90001  V
** inputVoltageBiasXXpXX2: 4.28101  V
** out: 2.5  V
** outFirstStage: 4.26401  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.62801  V
** innerTransistorStack1Load2: 4.62001  V
** innerTransistorStack2Load2: 4.62001  V
** out1: 4.26101  V
** sourceGCC1: 0.518001  V
** sourceGCC2: 0.518001  V
** sourceTransconductance: 3.27501  V
** innerStageBias: 0.635001  V


.END