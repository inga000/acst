** Name: one_stage_single_output_op_amp76

.MACRO one_stage_single_output_op_amp76 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=87e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=37e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=22e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=87e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=132e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=132e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=37e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageLoad12 out outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=235e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=336e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=305e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=305e-6
mFoldedCascodeFirstStageLoad16 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=336e-6
mMainBias17 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=38e-6
mMainBias18 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp76

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 3.55301 mW
** Area: 4486 (mu_m)^2
** Transit frequency: 8.48601 MHz
** Transit frequency with error factor: 8.48582 MHz
** Slew rate: 10.242 V/mu_s
** Phase margin: 87.6626°
** CMRR: 144 dB
** VoutMax: 4.01001 V
** VoutMin: 0.430001 V
** VcmMax: 5.17001 V
** VcmMin: 1.73001 V


** Expected Currents: 
** NormalTransistorPmos: -3.84409e+07 muA
** NormalTransistorPmos: -3.37959e+07 muA
** NormalTransistorPmos: -2.06154e+08 muA
** NormalTransistorPmos: -3.0923e+08 muA
** NormalTransistorPmos: -2.06155e+08 muA
** NormalTransistorPmos: -3.09231e+08 muA
** DiodeTransistorNmos: 2.06155e+08 muA
** NormalTransistorNmos: 2.06156e+08 muA
** NormalTransistorNmos: 2.06155e+08 muA
** NormalTransistorNmos: 2.06154e+08 muA
** DiodeTransistorNmos: 2.06153e+08 muA
** NormalTransistorNmos: 1.03078e+08 muA
** NormalTransistorNmos: 1.03078e+08 muA
** DiodeTransistorNmos: 3.84411e+07 muA
** NormalTransistorNmos: 3.84411e+07 muA
** DiodeTransistorNmos: 3.37961e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outInputVoltageBiasXXnXX1: 1.53401  V
** outSourceVoltageBiasXXnXX1: 0.767001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 1.04001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.367001  V
** out1: 0.572001  V
** sourceGCC1: 4.22401  V
** sourceGCC2: 4.22401  V
** sourceTransconductance: 1.90201  V
** inner: 0.767001  V


.END