** Name: two_stage_single_output_op_amp_74_8

.MACRO two_stage_single_output_op_amp_74_8 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=161e-6
m2 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=93e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=43e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=57e-6
m5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
m6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=19e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=26e-6
m8 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=424e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=9e-6 W=95e-6
m10 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
m11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=12e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=12e-6
m13 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=43e-6
m14 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=511e-6
m15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=161e-6
m16 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=427e-6
m17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=186e-6
m18 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=296e-6
m19 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=414e-6
m20 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=186e-6
m21 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=105e-6
m22 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=105e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6e-12
.EOM two_stage_single_output_op_amp_74_8

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 9.10101 mW
** Area: 11546 (mu_m)^2
** Transit frequency: 4.65901 MHz
** Transit frequency with error factor: 4.65915 MHz
** Slew rate: 4.14352 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 1.07001 V
** VcmMax: 5.15001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorPmos: -1.14523e+08 muA
** NormalTransistorPmos: -1.59013e+08 muA
** NormalTransistorPmos: -2.51799e+07 muA
** NormalTransistorPmos: -4.07589e+07 muA
** NormalTransistorPmos: -2.51799e+07 muA
** NormalTransistorPmos: -4.07589e+07 muA
** NormalTransistorNmos: 2.51791e+07 muA
** NormalTransistorNmos: 2.51791e+07 muA
** DiodeTransistorNmos: 2.51791e+07 muA
** NormalTransistorNmos: 3.11551e+07 muA
** DiodeTransistorNmos: 3.11541e+07 muA
** NormalTransistorNmos: 1.55781e+07 muA
** NormalTransistorNmos: 1.55781e+07 muA
** NormalTransistorNmos: 1.44517e+09 muA
** NormalTransistorNmos: 1.44517e+09 muA
** NormalTransistorPmos: -1.44516e+09 muA
** DiodeTransistorNmos: 1.14524e+08 muA
** NormalTransistorNmos: 1.14525e+08 muA
** DiodeTransistorNmos: 1.59014e+08 muA
** DiodeTransistorNmos: 1.59015e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.22201  V
** outInputVoltageBiasXXnXX2: 1.37101  V
** outSourceVoltageBiasXXnXX1: 0.611001  V
** outSourceVoltageBiasXXnXX2: 0.721001  V
** outSourceVoltageBiasXXpXX1: 4.18201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.611001  V
** out1: 1.18401  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.91901  V
** innerStageBias: 0.617001  V
** inner: 0.612001  V


.END