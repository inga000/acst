** Name: two_stage_single_output_op_amp_147_7

.MACRO two_stage_single_output_op_amp_147_7 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=14e-6
m2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
m3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=12e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=8e-6
m5 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
m6 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=12e-6
m7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=28e-6
m8 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=25e-6
m9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
m10 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=28e-6
m11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=75e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=412e-6
m13 outFirstStage outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=74e-6
m14 FirstStageYinnerOutputLoad1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=74e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 11.2001e-12
.EOM two_stage_single_output_op_amp_147_7

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 3.91901 mW
** Area: 4040 (mu_m)^2
** Transit frequency: 5.03901 MHz
** Transit frequency with error factor: 5.01796 MHz
** Slew rate: 4.74935 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.76001 V
** VoutMin: 0.180001 V
** VcmMax: 4.79001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorNmos: 1.78961e+07 muA
** DiodeTransistorNmos: 1.36574e+08 muA
** DiodeTransistorNmos: 1.36574e+08 muA
** NormalTransistorNmos: 1.36574e+08 muA
** NormalTransistorNmos: 1.36574e+08 muA
** NormalTransistorPmos: -1.63238e+08 muA
** NormalTransistorPmos: -1.63238e+08 muA
** NormalTransistorNmos: 5.33291e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 4.29522e+08 muA
** NormalTransistorPmos: -4.29521e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.78969e+07 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.19401  V
** outVoltageBiasXXpXX1: 3.82501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.28401  V
** innerSourceLoad1: 1.14201  V
** innerTransistorStack2Load1: 1.14201  V
** sourceTransconductance: 1.94501  V


.END