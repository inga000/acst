** Name: two_stage_single_output_op_amp_72_7

.MACRO two_stage_single_output_op_amp_72_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=76e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=64e-6
mFoldedCascodeFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=40e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=48e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=13e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=13e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=40e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=64e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=185e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=76e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=19e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=114e-6
mFoldedCascodeFirstStageLoad17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=19e-6
mMainBias18 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=306e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_72_7

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 7.93801 mW
** Area: 4312 (mu_m)^2
** Transit frequency: 5.95001 MHz
** Transit frequency with error factor: 5.94488 MHz
** Slew rate: 4.08418 V/mu_s
** Phase margin: 64.1713°
** CMRR: 109 dB
** VoutMax: 4.25 V
** VoutMin: 0.720001 V
** VcmMax: 5.17001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorPmos: -4.15689e+07 muA
** NormalTransistorPmos: -3.05639e+08 muA
** NormalTransistorPmos: -1.84589e+07 muA
** NormalTransistorPmos: -3.14299e+07 muA
** NormalTransistorPmos: -1.84589e+07 muA
** NormalTransistorPmos: -3.14299e+07 muA
** DiodeTransistorNmos: 1.84581e+07 muA
** NormalTransistorNmos: 1.84581e+07 muA
** NormalTransistorNmos: 2.59391e+07 muA
** DiodeTransistorNmos: 2.59381e+07 muA
** NormalTransistorNmos: 1.29701e+07 muA
** NormalTransistorNmos: 1.29701e+07 muA
** NormalTransistorNmos: 1.15749e+09 muA
** NormalTransistorPmos: -1.15748e+09 muA
** DiodeTransistorNmos: 4.15681e+07 muA
** NormalTransistorNmos: 4.15671e+07 muA
** DiodeTransistorNmos: 3.0564e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.16001  V
** outSourceVoltageBiasXXnXX1: 0.580001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 1.12701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.556001  V
** sourceGCC1: 4.19401  V
** sourceGCC2: 4.19401  V
** sourceTransconductance: 1.94101  V
** inner: 0.579001  V


.END