** Name: symmetrical_op_amp154

.MACRO symmetrical_op_amp154 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=9e-6
mMainBias2 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=24e-6
mSecondStage1StageBias3 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=94e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=6e-6 W=94e-6
mSymmetricalFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=78e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=43e-6
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=43e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=120e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=5e-6 W=120e-6
mSymmetricalFirstStageLoad10 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=51e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=123e-6
mSecondStage1Transconductor12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=123e-6
mSymmetricalFirstStageLoad13 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=51e-6
mSymmetricalFirstStageStageBias14 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=78e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias15 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=94e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=24e-6
mSymmetricalFirstStageTransconductor17 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=23e-6
mSecondStage1StageBias18 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=6e-6 W=94e-6
mSymmetricalFirstStageTransconductor19 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=23e-6
mMainBias20 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=30e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp154

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 0.784001 mW
** Area: 6822 (mu_m)^2
** Transit frequency: 2.57801 MHz
** Transit frequency with error factor: 2.5784 MHz
** Slew rate: 4.56005 V/mu_s
** Phase margin: 70.4739°
** CMRR: 144 dB
** negPSRR: 49 dB
** posPSRR: 70 dB
** VoutMax: 3.62001 V
** VoutMin: 0.310001 V
** VcmMax: 3.06001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.24859e+07 muA
** NormalTransistorNmos: 1.64781e+07 muA
** NormalTransistorNmos: 1.64771e+07 muA
** NormalTransistorNmos: 1.64781e+07 muA
** NormalTransistorNmos: 1.64771e+07 muA
** NormalTransistorPmos: -3.29579e+07 muA
** DiodeTransistorPmos: -3.29569e+07 muA
** NormalTransistorPmos: -1.64789e+07 muA
** NormalTransistorPmos: -1.64789e+07 muA
** NormalTransistorNmos: 4.57111e+07 muA
** NormalTransistorNmos: 4.57121e+07 muA
** NormalTransistorPmos: -4.57119e+07 muA
** DiodeTransistorPmos: -4.57129e+07 muA
** DiodeTransistorPmos: -4.57119e+07 muA
** NormalTransistorPmos: -4.57129e+07 muA
** NormalTransistorNmos: 4.57111e+07 muA
** NormalTransistorNmos: 4.57121e+07 muA
** DiodeTransistorNmos: 1.24851e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.34001  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 4.03001  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 3.06001  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.717001  V
** outSourceVoltageBiasXXpXX1: 4.17101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.160001  V
** innerTransistorStack2Load1: 0.160001  V
** sourceTransconductance: 3.34601  V
** innerTransconductance: 0.150001  V
** inner: 4.02701  V
** inner: 0.150001  V
** inner: 4.16801  V


.END