.suckt  two_stage_single_output_op_amp_143_7 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
m3 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos
m5 FirstStageYout1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m6 outFirstStage inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c2 out sourceNmos 
m10 out ibias sourceNmos sourceNmos nmos
m11 out outFirstStage sourcePmos sourcePmos pmos
m12 ibias ibias sourceNmos sourceNmos nmos
m13 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_143_7

