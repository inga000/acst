.suckt  two_stage_single_output_op_amp_107_10 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mMainBias2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mMainBias3 outVoltageBiasXXpXX3 ibias sourceNmos sourceNmos nmos
mMainBias4 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mTelescopicFirstStageLoad5 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mTelescopicFirstStageLoad6 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mTelescopicFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
mTelescopicFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos
mTelescopicFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mTelescopicFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos
mTelescopicFirstStageStageBias11 sourceTransconductance outVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
mTelescopicFirstStageStageBias12 FirstStageYinnerStageBias outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias15 out ibias sourceNmos sourceNmos nmos
mSecondStage1Transconductor16 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
mMainBias18 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias19 ibias ibias sourceNmos sourceNmos nmos
mMainBias20 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
mSecondStage1StageBias21 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mMainBias22 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_107_10

