** Name: two_stage_single_output_op_amp_60_8

.MACRO two_stage_single_output_op_amp_60_8 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=40e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=45e-6
m3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=21e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=84e-6
m5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=408e-6
m6 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=347e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=14e-6
m8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=14e-6
m9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=31e-6
m10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=31e-6
m11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=507e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=194e-6
m13 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=177e-6
m14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=6e-6 W=519e-6
m15 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=408e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=140e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=140e-6
m18 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=84e-6
m19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_60_8

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 5.99601 mW
** Area: 12828 (mu_m)^2
** Transit frequency: 5.46201 MHz
** Transit frequency with error factor: 5.46211 MHz
** Slew rate: 8.30948 V/mu_s
** Phase margin: 63.5984°
** CMRR: 142 dB
** VoutMax: 4.25 V
** VoutMin: 0.740001 V
** VcmMax: 3.05001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -8.57089e+07 muA
** NormalTransistorNmos: 3.86611e+07 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorNmos: 3.86601e+07 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorPmos: -3.86619e+07 muA
** NormalTransistorPmos: -3.86609e+07 muA
** DiodeTransistorPmos: -3.86619e+07 muA
** NormalTransistorPmos: -4.07649e+07 muA
** DiodeTransistorPmos: -4.07639e+07 muA
** NormalTransistorPmos: -2.03829e+07 muA
** NormalTransistorPmos: -2.03829e+07 muA
** NormalTransistorNmos: 9.754e+08 muA
** NormalTransistorNmos: 9.75399e+08 muA
** NormalTransistorPmos: -9.75399e+08 muA
** DiodeTransistorNmos: 8.57081e+07 muA
** DiodeTransistorNmos: 8.57091e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.30201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11901  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.25701  V
** out1: 3.53501  V
** sourceGCC1: 0.533001  V
** sourceGCC2: 0.533001  V
** sourceTransconductance: 3.31901  V
** innerStageBias: 0.531001  V
** inner: 4.14801  V


.END