** Name: two_stage_single_output_op_amp_130_3

.MACRO two_stage_single_output_op_amp_130_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=7e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=9e-6 W=41e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=176e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=29e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=101e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=101e-6
mSimpleFirstStageLoad8 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=99e-6
mMainBias9 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=454e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=65e-6
mSimpleFirstStageLoad11 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=99e-6
mMainBias12 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=295e-6
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=53e-6
mSimpleFirstStageLoad14 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=9e-6 W=41e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=362e-6
mSecondStage1StageBias17 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=597e-6
mSimpleFirstStageLoad18 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=9e-6
mSimpleFirstStageTransconductor19 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=53e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_130_3

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 9.32001 mW
** Area: 5420 (mu_m)^2
** Transit frequency: 4.98901 MHz
** Transit frequency with error factor: 4.97931 MHz
** Slew rate: 23.6279 V/mu_s
** Phase margin: 73.9116°
** CMRR: 77 dB
** VoutMax: 4.33001 V
** VoutMin: 0.410001 V
** VcmMax: 3.31001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 2.94448e+08 muA
** NormalTransistorNmos: 4.49135e+08 muA
** NormalTransistorPmos: -4.56909e+07 muA
** NormalTransistorPmos: -4.56899e+07 muA
** DiodeTransistorPmos: -4.56909e+07 muA
** NormalTransistorNmos: 9.95031e+07 muA
** NormalTransistorNmos: 9.95021e+07 muA
** NormalTransistorNmos: 9.95021e+07 muA
** NormalTransistorNmos: 9.95021e+07 muA
** NormalTransistorPmos: -1.07626e+08 muA
** NormalTransistorPmos: -5.38129e+07 muA
** NormalTransistorPmos: -5.38129e+07 muA
** NormalTransistorNmos: 9.1131e+08 muA
** NormalTransistorPmos: -9.11309e+08 muA
** NormalTransistorPmos: -9.1131e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.94447e+08 muA
** DiodeTransistorPmos: -4.49134e+08 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.06001  V
** out: 2.5  V
** outFirstStage: 0.814001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.587001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.587001  V
** out1: 2.37201  V
** sourceTransconductance: 3.81401  V
** innerStageBias: 4.54101  V


.END