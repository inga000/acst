** Name: two_stage_single_output_op_amp_33_10

.MACRO two_stage_single_output_op_amp_33_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=58e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=365e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=87e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=76e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=17e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=39e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=9e-6 W=291e-6
mMainBias9 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=267e-6
mSecondStage1StageBias10 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=532e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=17e-6
mMainBias12 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=365e-6
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=399e-6
mSecondStage1Transconductor15 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=600e-6
mSimpleFirstStageLoad16 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=72e-6
mMainBias17 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=334e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.60001e-12
.EOM two_stage_single_output_op_amp_33_10

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 7.46601 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 7.13801 MHz
** Transit frequency with error factor: 7.13443 MHz
** Slew rate: 6.72724 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** negPSRR: 105 dB
** posPSRR: 100 dB
** VoutMax: 4.25 V
** VoutMin: 0.240001 V
** VcmMax: 4.46001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 1.96341e+07 muA
** NormalTransistorNmos: 4.41673e+08 muA
** NormalTransistorPmos: -8.64109e+07 muA
** DiodeTransistorPmos: -3.23799e+07 muA
** NormalTransistorPmos: -3.23799e+07 muA
** NormalTransistorPmos: -3.23799e+07 muA
** NormalTransistorNmos: 6.47571e+07 muA
** NormalTransistorNmos: 6.47561e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 8.70761e+08 muA
** NormalTransistorPmos: -8.7076e+08 muA
** NormalTransistorPmos: -8.70761e+08 muA
** DiodeTransistorNmos: 8.64101e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.96349e+07 muA
** DiodeTransistorPmos: -4.41672e+08 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.08701  V
** outVoltageBiasXXnXX1: 0.801001  V
** outVoltageBiasXXpXX0: 4.07401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.27801  V
** innerStageBias: 0.242001  V
** innerTransistorStack2Load1: 4.47401  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.65101  V


.END