** Name: two_stage_single_output_op_amp_75_1

.MACRO two_stage_single_output_op_amp_75_1 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=22e-6
m2 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=14e-6
m3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=76e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=29e-6
m5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=29e-6
m6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=180e-6
m7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=22e-6
m8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=340e-6
m9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=340e-6
m10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=72e-6
m11 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
m12 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=140e-6
m13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=411e-6
m14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=108e-6
m15 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=322e-6
m16 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=74e-6
m17 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=74e-6
m18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=559e-6
m19 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=322e-6
m20 outVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=190e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 13.3001e-12
.EOM two_stage_single_output_op_amp_75_1

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 13.7341 mW
** Area: 14998 (mu_m)^2
** Transit frequency: 10.2451 MHz
** Transit frequency with error factor: 10.2446 MHz
** Slew rate: 9.65531 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 4.62001 V
** VoutMin: 0.340001 V
** VcmMax: 5.02001 V
** VcmMin: 1.5 V


** Expected Currents: 
** NormalTransistorNmos: 2.94448e+08 muA
** NormalTransistorNmos: 7.75891e+07 muA
** NormalTransistorPmos: -5.0835e+08 muA
** NormalTransistorPmos: -1.29516e+08 muA
** NormalTransistorPmos: -1.94273e+08 muA
** NormalTransistorPmos: -1.29519e+08 muA
** NormalTransistorPmos: -1.94278e+08 muA
** DiodeTransistorNmos: 1.29519e+08 muA
** NormalTransistorNmos: 1.2952e+08 muA
** NormalTransistorNmos: 1.29519e+08 muA
** NormalTransistorNmos: 1.29516e+08 muA
** NormalTransistorNmos: 1.29515e+08 muA
** NormalTransistorNmos: 6.47581e+07 muA
** NormalTransistorNmos: 6.47581e+07 muA
** NormalTransistorNmos: 1.46785e+09 muA
** NormalTransistorPmos: -1.46784e+09 muA
** DiodeTransistorNmos: 5.08351e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.94447e+08 muA
** DiodeTransistorPmos: -7.75899e+07 muA


** Expected Voltages: 
** ibias: 0.564001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.744001  V
** outVoltageBiasXXnXX1: 1.14801  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.05101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.359001  V
** innerTransistorStack2Load2: 0.466001  V
** out1: 0.668001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V


.END