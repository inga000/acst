** Name: two_stage_single_output_op_amp_197_7

.MACRO two_stage_single_output_op_amp_197_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=20e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=54e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=11e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=48e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=22e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=391e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=20e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=48e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=176e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=176e-6
mSimpleFirstStageLoad16 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=455e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=395e-6
mSimpleFirstStageLoad18 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=455e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=50e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=9e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_197_7

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 5.99301 mW
** Area: 11863 (mu_m)^2
** Transit frequency: 4.62701 MHz
** Transit frequency with error factor: 4.62328 MHz
** Slew rate: 4.36049 V/mu_s
** Phase margin: 60.1606°
** CMRR: 120 dB
** VoutMax: 4.25 V
** VoutMin: 0.310001 V
** VcmMax: 4.59001 V
** VcmMin: 1.55001 V


** Expected Currents: 
** NormalTransistorPmos: -4.62149e+07 muA
** NormalTransistorPmos: -8.15499e+06 muA
** DiodeTransistorNmos: 1.50863e+08 muA
** DiodeTransistorNmos: 1.50862e+08 muA
** NormalTransistorNmos: 1.50861e+08 muA
** NormalTransistorNmos: 1.50862e+08 muA
** NormalTransistorPmos: -1.61021e+08 muA
** NormalTransistorPmos: -1.6102e+08 muA
** NormalTransistorPmos: -1.61019e+08 muA
** NormalTransistorPmos: -1.6102e+08 muA
** NormalTransistorNmos: 2.03171e+07 muA
** NormalTransistorNmos: 2.03161e+07 muA
** NormalTransistorNmos: 1.01591e+07 muA
** NormalTransistorNmos: 1.01591e+07 muA
** NormalTransistorNmos: 8.02119e+08 muA
** NormalTransistorPmos: -8.02118e+08 muA
** DiodeTransistorNmos: 4.62141e+07 muA
** DiodeTransistorNmos: 8.15401e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 3.93001  V
** outVoltageBiasXXnXX1: 1.09301  V
** outVoltageBiasXXnXX2: 0.715001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.14901  V
** innerStageBias: 0.411001  V
** innerTransistorStack1Load2: 4.01601  V
** innerTransistorStack2Load1: 1.15001  V
** innerTransistorStack2Load2: 4.01601  V
** out1: 2.15401  V
** sourceTransconductance: 1.94501  V


.END