** Name: two_stage_single_output_op_amp_57_12

.MACRO two_stage_single_output_op_amp_57_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=15e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=10e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=336e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=38e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=10e-6 W=36e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=45e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=45e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=15e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=336e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=10e-6 W=36e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=24e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=599e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=158e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=158e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=394e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mMainBias20 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=228e-6
mMainBias21 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=157e-6
mSecondStage1Transconductor22 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=484e-6
mFoldedCascodeFirstStageLoad23 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.6001e-12
.EOM two_stage_single_output_op_amp_57_12

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 9.85101 mW
** Area: 14996 (mu_m)^2
** Transit frequency: 6.40501 MHz
** Transit frequency with error factor: 6.39839 MHz
** Slew rate: 8.2035 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** VoutMax: 4.25 V
** VoutMin: 1.71001 V
** VcmMax: 3.19001 V
** VcmMin: 0.140001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -6.07539e+07 muA
** NormalTransistorPmos: -4.17749e+07 muA
** NormalTransistorNmos: 1.1173e+08 muA
** NormalTransistorNmos: 1.91538e+08 muA
** NormalTransistorNmos: 1.11728e+08 muA
** NormalTransistorNmos: 1.91534e+08 muA
** DiodeTransistorPmos: -1.11727e+08 muA
** NormalTransistorPmos: -1.11727e+08 muA
** NormalTransistorPmos: -1.59613e+08 muA
** NormalTransistorPmos: -1.59612e+08 muA
** NormalTransistorPmos: -7.98069e+07 muA
** NormalTransistorPmos: -7.98069e+07 muA
** NormalTransistorNmos: 1.36311e+09 muA
** DiodeTransistorNmos: 1.36311e+09 muA
** NormalTransistorPmos: -1.3631e+09 muA
** NormalTransistorPmos: -1.3631e+09 muA
** DiodeTransistorNmos: 6.07531e+07 muA
** NormalTransistorNmos: 6.07521e+07 muA
** DiodeTransistorNmos: 4.17741e+07 muA
** DiodeTransistorNmos: 4.17751e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.11801  V
** inputVoltageBiasXXnXX2: 2.21501  V
** out: 2.5  V
** outFirstStage: 4.08101  V
** outSourceVoltageBiasXXnXX1: 1.05901  V
** outSourceVoltageBiasXXnXX2: 1.11101  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40001  V
** out1: 4.07001  V
** sourceGCC1: 1.20201  V
** sourceGCC2: 1.20201  V
** sourceTransconductance: 3.35401  V
** innerTransconductance: 4.64501  V
** inner: 1.05401  V


.END