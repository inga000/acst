** Name: two_stage_single_output_op_amp_151_9

.MACRO two_stage_single_output_op_amp_151_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=6e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=5e-6 W=6e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=24e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=266e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=200e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=6e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=54e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=24e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=266e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=6e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=54e-6
mSimpleFirstStageLoad14 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=74e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=147e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=596e-6
mSimpleFirstStageLoad17 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=74e-6
mMainBias18 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=228e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.40001e-12
.EOM two_stage_single_output_op_amp_151_9

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 10.0701 mW
** Area: 8684 (mu_m)^2
** Transit frequency: 6.78601 MHz
** Transit frequency with error factor: 6.7688 MHz
** Slew rate: 6.3955 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 1.86001 V
** VcmMax: 5.18001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorPmos: -1.35525e+08 muA
** NormalTransistorPmos: -2.10203e+08 muA
** DiodeTransistorNmos: 4.71421e+07 muA
** NormalTransistorNmos: 4.71411e+07 muA
** NormalTransistorNmos: 4.71421e+07 muA
** DiodeTransistorNmos: 4.71411e+07 muA
** NormalTransistorPmos: -6.77129e+07 muA
** NormalTransistorPmos: -6.77129e+07 muA
** NormalTransistorNmos: 4.11391e+07 muA
** NormalTransistorNmos: 2.05701e+07 muA
** NormalTransistorNmos: 2.05701e+07 muA
** NormalTransistorNmos: 1.51286e+09 muA
** DiodeTransistorNmos: 1.51286e+09 muA
** NormalTransistorPmos: -1.51285e+09 muA
** DiodeTransistorNmos: 1.35526e+08 muA
** NormalTransistorNmos: 1.35525e+08 muA
** DiodeTransistorNmos: 2.10204e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.27001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 1.13501  V
** outVoltageBiasXXnXX2: 0.563001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.01201  V
** innerTransistorStack1Load1: 1.00601  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 1.13101  V


.END