** Name: symmetrical_op_amp80

.MACRO symmetrical_op_amp80 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=20e-6
m2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
m3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=3e-6 W=208e-6
m4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
m5 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m6 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=117e-6
m7 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=117e-6
m8 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=200e-6
m9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=47e-6
m10 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=159e-6
m11 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=47e-6
m12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=600e-6
m13 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=20e-6
m15 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=599e-6
m16 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
m17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=265e-6
m18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=265e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp80

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 5.43901 mW
** Area: 9167 (mu_m)^2
** Transit frequency: 27.4451 MHz
** Transit frequency with error factor: 27.4448 MHz
** Slew rate: 33.816 V/mu_s
** Phase margin: 65.8902°
** CMRR: 146 dB
** negPSRR: 62 dB
** posPSRR: 55 dB
** VoutMax: 4.56001 V
** VoutMin: 1.23001 V
** VcmMax: 4.57001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 9.95911e+07 muA
** DiodeTransistorPmos: -1.48151e+08 muA
** DiodeTransistorPmos: -1.48151e+08 muA
** NormalTransistorNmos: 2.96302e+08 muA
** DiodeTransistorNmos: 2.96301e+08 muA
** NormalTransistorNmos: 1.48152e+08 muA
** NormalTransistorNmos: 1.48152e+08 muA
** NormalTransistorNmos: 3.41003e+08 muA
** NormalTransistorNmos: 3.41002e+08 muA
** NormalTransistorPmos: -3.41002e+08 muA
** NormalTransistorPmos: -3.41001e+08 muA
** DiodeTransistorNmos: 3.41001e+08 muA
** DiodeTransistorNmos: 3.41e+08 muA
** NormalTransistorPmos: -3.41e+08 muA
** NormalTransistorPmos: -3.41001e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.95919e+07 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceStageBiasComplementarySecondStage: 0.952001  V
** inSourceTransconductanceComplementarySecondStage: 4.16901  V
** innerComplementarySecondStage: 1.59701  V
** out: 2.5  V
** outFirstStage: 4.16901  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.90201  V
** innerStageBias: 0.915001  V
** innerTransconductance: 4.42801  V
** inner: 4.42801  V
** inner: 0.556001  V


.END