** Name: two_stage_single_output_op_amp_137_5

.MACRO two_stage_single_output_op_amp_137_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=10e-6 W=127e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=127e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=113e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=312e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=128e-6
mSimpleFirstStageLoad7 FirstStageYout1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=503e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=471e-6
mSimpleFirstStageLoad9 outFirstStage ibias sourceNmos sourceNmos nmos4 L=2e-6 W=503e-6
mMainBias10 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=295e-6
mMainBias11 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=231e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=10e-6 W=127e-6
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=306e-6
mSimpleFirstStageStageBias14 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=449e-6
mMainBias15 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=113e-6
mSecondStage1StageBias16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=312e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=127e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=306e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.3001e-12
.EOM two_stage_single_output_op_amp_137_5

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 12.9771 mW
** Area: 14912 (mu_m)^2
** Transit frequency: 11.3181 MHz
** Transit frequency with error factor: 11.2634 MHz
** Slew rate: 24.5923 V/mu_s
** Phase margin: 60.1606°
** CMRR: 71 dB
** VoutMax: 3.04001 V
** VoutMin: 0.150001 V
** VcmMax: 3.11001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorNmos: 3.24691e+08 muA
** NormalTransistorNmos: 2.57296e+08 muA
** DiodeTransistorPmos: -1.09342e+08 muA
** NormalTransistorPmos: -1.09343e+08 muA
** NormalTransistorPmos: -1.09342e+08 muA
** DiodeTransistorPmos: -1.09343e+08 muA
** NormalTransistorNmos: 5.53191e+08 muA
** NormalTransistorNmos: 5.53191e+08 muA
** NormalTransistorPmos: -8.87696e+08 muA
** NormalTransistorPmos: -4.43847e+08 muA
** NormalTransistorPmos: -4.43847e+08 muA
** NormalTransistorNmos: 8.9708e+08 muA
** NormalTransistorPmos: -8.97079e+08 muA
** DiodeTransistorPmos: -8.9708e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.2469e+08 muA
** NormalTransistorPmos: -3.24691e+08 muA
** DiodeTransistorPmos: -2.57295e+08 muA


** Expected Voltages: 
** ibias: 0.567001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.47601  V
** outSourceVoltageBiasXXpXX1: 3.73801  V
** outVoltageBiasXXpXX2: 3.85801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.73901  V
** innerTransistorStack1Load1: 3.73801  V
** out1: 2.95501  V
** sourceTransconductance: 3.81401  V
** inner: 3.73201  V


.END