** Name: one_stage_single_output_op_amp75

.MACRO one_stage_single_output_op_amp75 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=97e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=39e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=6e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=23e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=139e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=97e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=75e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=75e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=100e-6
mFoldedCascodeFirstStageLoad11 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=93e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=121e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=105e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=105e-6
mMainBias15 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageLoad16 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=121e-6
mMainBias17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=49e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp75

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 1.51001 mW
** Area: 6097 (mu_m)^2
** Transit frequency: 2.66401 MHz
** Transit frequency with error factor: 2.66433 MHz
** Slew rate: 3.53985 V/mu_s
** Phase margin: 89.3815°
** CMRR: 139 dB
** VoutMax: 4.02001 V
** VoutMin: 0.490001 V
** VcmMax: 5.17001 V
** VcmMin: 1.46001 V


** Expected Currents: 
** NormalTransistorPmos: -4.88509e+07 muA
** NormalTransistorPmos: -2.02769e+07 muA
** NormalTransistorPmos: -7.09709e+07 muA
** NormalTransistorPmos: -1.06454e+08 muA
** NormalTransistorPmos: -7.09729e+07 muA
** NormalTransistorPmos: -1.06456e+08 muA
** DiodeTransistorNmos: 7.09711e+07 muA
** NormalTransistorNmos: 7.09721e+07 muA
** NormalTransistorNmos: 7.09711e+07 muA
** NormalTransistorNmos: 7.09691e+07 muA
** NormalTransistorNmos: 7.09681e+07 muA
** NormalTransistorNmos: 3.54851e+07 muA
** NormalTransistorNmos: 3.54851e+07 muA
** DiodeTransistorNmos: 4.88501e+07 muA
** DiodeTransistorNmos: 2.02761e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.639001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.09501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.485001  V
** innerTransistorStack2Load2: 0.478001  V
** out1: 0.683001  V
** sourceGCC1: 4.22401  V
** sourceGCC2: 4.22401  V
** sourceTransconductance: 1.88301  V


.END