** Name: two_stage_single_output_op_amp_108_7

.MACRO two_stage_single_output_op_amp_108_7 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=423e-6
m2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=105e-6
m3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=11e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=462e-6
m5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=110e-6
m6 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=479e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=109e-6
m8 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=128e-6
m9 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=109e-6
m10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=85e-6
m11 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=85e-6
m12 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=387e-6
m13 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=337e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=118e-6
m15 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=59e-6
m16 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=462e-6
m17 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=59e-6
m18 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=16e-6
m19 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=16e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 7.10001e-12
.EOM two_stage_single_output_op_amp_108_7

** Expected Performance Values: 
** Gain: 117 dB
** Power consumption: 12.6471 mW
** Area: 11281 (mu_m)^2
** Transit frequency: 2.56801 MHz
** Transit frequency with error factor: 2.56801 MHz
** Slew rate: 52.1525 V/mu_s
** Phase margin: 60.1606°
** CMRR: 126 dB
** VoutMax: 3 V
** VoutMin: 0.260001 V
** VcmMax: 3.02001 V
** VcmMin: -0.199999 V


** Expected Currents: 
** NormalTransistorNmos: 3.79499e+08 muA
** NormalTransistorPmos: -3.56792e+08 muA
** NormalTransistorPmos: -3.06672e+08 muA
** NormalTransistorPmos: -2.32189e+07 muA
** NormalTransistorPmos: -2.32189e+07 muA
** NormalTransistorNmos: 2.32181e+07 muA
** NormalTransistorNmos: 2.32171e+07 muA
** NormalTransistorNmos: 2.32181e+07 muA
** NormalTransistorNmos: 2.32171e+07 muA
** NormalTransistorPmos: -4.25939e+08 muA
** DiodeTransistorPmos: -4.25938e+08 muA
** NormalTransistorPmos: -2.32199e+07 muA
** NormalTransistorPmos: -2.32199e+07 muA
** NormalTransistorNmos: 1.41998e+09 muA
** NormalTransistorPmos: -1.41997e+09 muA
** DiodeTransistorNmos: 3.56793e+08 muA
** DiodeTransistorNmos: 3.06673e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -3.79498e+08 muA


** Expected Voltages: 
** ibias: 3.41801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXnXX2: 0.669001  V
** out: 2.5  V
** outFirstStage: 2.43601  V
** outSourceVoltageBiasXXpXX1: 4.21001  V
** outVoltageBiasXXpXX2: 2.27701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.46501  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 3.05001  V
** sourceGCC2: 3.05001  V
** inner: 4.20701  V


.END