.suckt  symmetrical_op_amp172 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m3 out2FirstStage out2FirstStage out1FirstStage out1FirstStage pmos
m4 out1FirstStage out1FirstStage sourcePmos sourcePmos pmos
m5 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage pmos
m6 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m7 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m8 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m9 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m10 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m11 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m12 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
m13 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m14 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m15 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos
m16 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos
m17 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m19 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m20 ibias ibias sourceNmos sourceNmos nmos
m21 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end symmetrical_op_amp172

