** Name: two_stage_single_output_op_amp_3_6

.MACRO two_stage_single_output_op_amp_3_6 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=89e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=20e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=231e-6
m7 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=599e-6
m8 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=339e-6
m9 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=207e-6
m10 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=89e-6
m11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
m12 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=231e-6
m13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=510e-6
m14 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
m15 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=108e-6
m16 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=510e-6
m17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
m18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.40001e-12
.EOM two_stage_single_output_op_amp_3_6

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 14.9461 mW
** Area: 14181 (mu_m)^2
** Transit frequency: 28.2121 MHz
** Transit frequency with error factor: 28.1631 MHz
** Slew rate: 77.0977 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** negPSRR: 90 dB
** posPSRR: 95 dB
** VoutMax: 3.02001 V
** VoutMin: 0.550001 V
** VcmMax: 3.68001 V
** VcmMin: 0.220001 V


** Expected Currents: 
** NormalTransistorNmos: 1.80961e+08 muA
** NormalTransistorPmos: -2.02769e+07 muA
** NormalTransistorPmos: -1.09497e+08 muA
** DiodeTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorNmos: 2.05013e+09 muA
** NormalTransistorNmos: 2.05013e+09 muA
** NormalTransistorPmos: -2.05012e+09 muA
** DiodeTransistorPmos: -2.05012e+09 muA
** DiodeTransistorNmos: 2.02761e+07 muA
** DiodeTransistorNmos: 1.09498e+08 muA
** DiodeTransistorPmos: -1.8096e+08 muA
** NormalTransistorPmos: -1.8096e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.605001  V
** outInputVoltageBiasXXpXX1: 2.45601  V
** outSourceVoltageBiasXXpXX1: 3.72801  V
** outVoltageBiasXXnXX0: 0.633001  V
** outVoltageBiasXXnXX1: 0.952001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 0.368001  V
** out1: 0.605001  V
** sourceTransconductance: 3.57901  V
** innerTransconductance: 0.200001  V
** inner: 3.72801  V


.END