** Name: two_stage_single_output_op_amp_151_8

.MACRO two_stage_single_output_op_amp_151_8 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=8e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
m6 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=372e-6
m7 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=8e-6
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=132e-6
m9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=132e-6
m11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
m12 SecondStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=593e-6
m13 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=245e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=434e-6
m15 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=163e-6
m16 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
m17 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=163e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10e-12
.EOM two_stage_single_output_op_amp_151_8

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 13.6751 mW
** Area: 6058 (mu_m)^2
** Transit frequency: 6.62001 MHz
** Transit frequency with error factor: 6.61053 MHz
** Slew rate: 6.23926 V/mu_s
** Phase margin: 60.1606°
** CMRR: 88 dB
** VoutMax: 4.25 V
** VoutMin: 0.560001 V
** VcmMax: 5.25 V
** VcmMin: 0.850001 V


** Expected Currents: 
** NormalTransistorPmos: -2.63565e+08 muA
** NormalTransistorPmos: -1.0576e+08 muA
** DiodeTransistorNmos: 3.97871e+07 muA
** NormalTransistorNmos: 3.97881e+07 muA
** NormalTransistorNmos: 3.97871e+07 muA
** DiodeTransistorNmos: 3.97881e+07 muA
** NormalTransistorPmos: -7.12149e+07 muA
** NormalTransistorPmos: -7.12149e+07 muA
** NormalTransistorNmos: 6.28531e+07 muA
** NormalTransistorNmos: 3.14271e+07 muA
** NormalTransistorNmos: 3.14271e+07 muA
** NormalTransistorNmos: 2.20329e+09 muA
** NormalTransistorNmos: 2.20329e+09 muA
** NormalTransistorPmos: -2.20328e+09 muA
** DiodeTransistorNmos: 2.63566e+08 muA
** DiodeTransistorNmos: 1.05761e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.700001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 0.964001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 1.09401  V
** innerTransistorStack2Load1: 1.09401  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.295001  V


.END