.suckt  one_stage_fully_differential_op_amp49 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m3 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m4 outFeedback outFeedback sourcePmos sourcePmos pmos
m5 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m6 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m7 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m8 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m9 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m10 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m11 out1 outFeedback sourcePmos sourcePmos pmos
m12 out2 outFeedback sourcePmos sourcePmos pmos
m13 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m14 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m15 out1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m16 out2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out1 sourceNmos 
c2 out2 sourceNmos 
m17 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m18 ibias ibias sourceNmos sourceNmos nmos
m19 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end one_stage_fully_differential_op_amp49

