** Name: two_stage_single_output_op_amp_73_9

.MACRO two_stage_single_output_op_amp_73_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=9e-6 W=9e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=7e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=282e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
m5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=21e-6
m6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=24e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
m8 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=282e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=5e-6 W=6e-6
m10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=17e-6
m11 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=21e-6
m12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=22e-6
m13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=22e-6
m14 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=9e-6 W=53e-6
m15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
m16 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=249e-6
m17 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=32e-6
m18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=156e-6
m19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=64e-6
m20 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=156e-6
m21 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=74e-6
m22 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=74e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 5.20001e-12
.EOM two_stage_single_output_op_amp_73_9

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 7.01101 mW
** Area: 6359 (mu_m)^2
** Transit frequency: 4.5 MHz
** Transit frequency with error factor: 4.50031 MHz
** Slew rate: 4.02283 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 4.25 V
** VoutMin: 1.43001 V
** VcmMax: 5.12001 V
** VcmMin: 1.68001 V


** Expected Currents: 
** NormalTransistorPmos: -3.09149e+07 muA
** NormalTransistorPmos: -1.53989e+07 muA
** NormalTransistorPmos: -2.11189e+07 muA
** NormalTransistorPmos: -3.59109e+07 muA
** NormalTransistorPmos: -2.11189e+07 muA
** NormalTransistorPmos: -3.59109e+07 muA
** NormalTransistorNmos: 2.11181e+07 muA
** NormalTransistorNmos: 2.11181e+07 muA
** DiodeTransistorNmos: 2.11181e+07 muA
** NormalTransistorNmos: 2.95811e+07 muA
** NormalTransistorNmos: 2.95801e+07 muA
** NormalTransistorNmos: 1.47911e+07 muA
** NormalTransistorNmos: 1.47911e+07 muA
** NormalTransistorNmos: 1.2641e+09 muA
** DiodeTransistorNmos: 1.2641e+09 muA
** NormalTransistorPmos: -1.26409e+09 muA
** DiodeTransistorNmos: 3.09141e+07 muA
** NormalTransistorNmos: 3.09131e+07 muA
** DiodeTransistorNmos: 1.53981e+07 muA
** DiodeTransistorNmos: 1.53971e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.66301  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.83401  V
** outSourceVoltageBiasXXnXX1: 0.917001  V
** outSourceVoltageBiasXXnXX2: 0.833001  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.593001  V
** innerStageBias: 1.01401  V
** out1: 1.45201  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.89501  V
** inner: 0.916001  V


.END