** Name: two_stage_single_output_op_amp_206_8

.MACRO two_stage_single_output_op_amp_206_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=51e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=51e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=49e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=154e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=54e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=47e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=51e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=42e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=54e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=531e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=154e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=414e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=51e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=42e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=423e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=423e-6
mSimpleFirstStageLoad19 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=600e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=94e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=106e-6
mSimpleFirstStageLoad22 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=600e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=90e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.60001e-12
.EOM two_stage_single_output_op_amp_206_8

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 10.6361 mW
** Area: 8063 (mu_m)^2
** Transit frequency: 5.85301 MHz
** Transit frequency with error factor: 5.84861 MHz
** Slew rate: 5.51617 V/mu_s
** Phase margin: 60.1606°
** CMRR: 125 dB
** VoutMax: 4.25 V
** VoutMin: 0.730001 V
** VcmMax: 4.97001 V
** VcmMin: 1.43001 V


** Expected Currents: 
** NormalTransistorPmos: -8.98589e+07 muA
** NormalTransistorPmos: -9.34219e+07 muA
** DiodeTransistorNmos: 4.07813e+08 muA
** NormalTransistorNmos: 4.07814e+08 muA
** NormalTransistorNmos: 4.07815e+08 muA
** DiodeTransistorNmos: 4.07814e+08 muA
** NormalTransistorPmos: -4.23811e+08 muA
** NormalTransistorPmos: -4.23812e+08 muA
** NormalTransistorPmos: -4.23813e+08 muA
** NormalTransistorPmos: -4.23812e+08 muA
** NormalTransistorNmos: 3.19971e+07 muA
** DiodeTransistorNmos: 3.19961e+07 muA
** NormalTransistorNmos: 1.59991e+07 muA
** NormalTransistorNmos: 1.59991e+07 muA
** NormalTransistorNmos: 1.07627e+09 muA
** NormalTransistorNmos: 1.07626e+09 muA
** NormalTransistorPmos: -1.07626e+09 muA
** DiodeTransistorNmos: 8.98581e+07 muA
** NormalTransistorNmos: 8.98591e+07 muA
** DiodeTransistorNmos: 9.34211e+07 muA
** DiodeTransistorNmos: 9.34221e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.11401  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.28201  V
** outSourceVoltageBiasXXnXX1: 0.641001  V
** outSourceVoltageBiasXXnXX2: 0.559001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack1Load1: 1.15601  V
** innerTransistorStack1Load2: 4.16001  V
** innerTransistorStack2Load2: 4.16001  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.533001  V
** inner: 0.642001  V


.END