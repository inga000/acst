** Name: two_stage_single_output_op_amp_15_1

.MACRO two_stage_single_output_op_amp_15_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=28e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=61e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=9e-6
mMainBias5 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=190e-6
mSimpleFirstStageLoad7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=28e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=96e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=9e-6 W=38e-6
mSecondStage1StageBias11 out ibias sourcePmos sourcePmos pmos4 L=4e-6 W=564e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mMainBias13 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=14e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_15_1

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 0.710001 mW
** Area: 4619 (mu_m)^2
** Transit frequency: 2.65001 MHz
** Transit frequency with error factor: 2.64499 MHz
** Slew rate: 3.5001 V/mu_s
** Phase margin: 63.0254°
** CMRR: 98 dB
** negPSRR: 100 dB
** posPSRR: 173 dB
** VoutMax: 4.81001 V
** VoutMin: 0.150001 V
** VcmMax: 3.01001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 1.00131e+07 muA
** NormalTransistorPmos: -2.32799e+06 muA
** DiodeTransistorNmos: 7.89501e+06 muA
** NormalTransistorNmos: 7.89501e+06 muA
** NormalTransistorPmos: -1.57929e+07 muA
** NormalTransistorPmos: -1.57939e+07 muA
** NormalTransistorPmos: -7.89599e+06 muA
** NormalTransistorPmos: -7.89599e+06 muA
** NormalTransistorNmos: 9.38221e+07 muA
** NormalTransistorPmos: -9.38229e+07 muA
** DiodeTransistorNmos: 2.32701e+06 muA
** DiodeTransistorPmos: -1.00139e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.557001  V
** outVoltageBiasXXnXX0: 0.571001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.70601  V
** out1: 0.557001  V
** sourceTransconductance: 3.27401  V


.END