** Name: two_stage_single_output_op_amp_188_8

.MACRO two_stage_single_output_op_amp_188_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=10e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=22e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mSimpleFirstStageTransconductor7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=52e-6
mSimpleFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=18e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=291e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=545e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=5e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=52e-6
mSimpleFirstStageLoad15 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=102e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=425e-6
mSimpleFirstStageLoad17 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=102e-6
mMainBias18 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
mMainBias19 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_188_8

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 11.9321 mW
** Area: 3488 (mu_m)^2
** Transit frequency: 11.5771 MHz
** Transit frequency with error factor: 11.549 MHz
** Slew rate: 10.9115 V/mu_s
** Phase margin: 61.3065°
** CMRR: 91 dB
** VoutMax: 4.25 V
** VoutMin: 1.13001 V
** VcmMax: 5.21001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorPmos: -2.77049e+07 muA
** NormalTransistorPmos: -4.37239e+07 muA
** NormalTransistorNmos: 4.39621e+07 muA
** NormalTransistorNmos: 4.39631e+07 muA
** DiodeTransistorNmos: 4.39621e+07 muA
** NormalTransistorPmos: -6.87239e+07 muA
** NormalTransistorPmos: -6.87239e+07 muA
** NormalTransistorNmos: 4.95211e+07 muA
** DiodeTransistorNmos: 4.95201e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.1576e+09 muA
** NormalTransistorNmos: 2.1576e+09 muA
** NormalTransistorPmos: -2.15759e+09 muA
** DiodeTransistorNmos: 2.77041e+07 muA
** NormalTransistorNmos: 2.77031e+07 muA
** DiodeTransistorNmos: 4.37231e+07 muA
** DiodeTransistorNmos: 4.37221e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.17001  V
** outInputVoltageBiasXXnXX2: 1.44301  V
** outSourceVoltageBiasXXnXX1: 0.585001  V
** outSourceVoltageBiasXXnXX2: 0.822001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.12901  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.731001  V
** inner: 0.584001  V


.END