** Name: two_stage_single_output_op_amp_16_3

.MACRO two_stage_single_output_op_amp_16_3 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=39e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=30e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=21e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=203e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=33e-6
mMainBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=555e-6
mSimpleFirstStageLoad8 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=39e-6
mMainBias9 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=121e-6
mSimpleFirstStageTransconductor10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=33e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=370e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=203e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=595e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mMainBias16 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_16_3

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 2.66901 mW
** Area: 5014 (mu_m)^2
** Transit frequency: 2.64901 MHz
** Transit frequency with error factor: 2.64747 MHz
** Slew rate: 3.50007 V/mu_s
** Phase margin: 83.0789°
** CMRR: 98 dB
** negPSRR: 100 dB
** posPSRR: 172 dB
** VoutMax: 4.01001 V
** VoutMin: 0.150001 V
** VcmMax: 3.33001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 9.85511e+07 muA
** NormalTransistorPmos: -2.43329e+07 muA
** DiodeTransistorNmos: 7.90201e+06 muA
** NormalTransistorNmos: 7.90201e+06 muA
** NormalTransistorPmos: -1.58069e+07 muA
** DiodeTransistorPmos: -1.58079e+07 muA
** NormalTransistorPmos: -7.90299e+06 muA
** NormalTransistorPmos: -7.90299e+06 muA
** NormalTransistorNmos: 3.75136e+08 muA
** NormalTransistorPmos: -3.75135e+08 muA
** NormalTransistorPmos: -3.75134e+08 muA
** DiodeTransistorNmos: 2.43321e+07 muA
** DiodeTransistorPmos: -9.85519e+07 muA
** NormalTransistorPmos: -9.85529e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.559001  V
** outInputVoltageBiasXXpXX1: 3.54401  V
** outSourceVoltageBiasXXpXX1: 4.27201  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.664001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.559001  V
** sourceTransconductance: 3.27401  V
** innerStageBias: 4.22201  V
** inner: 4.27201  V


.END