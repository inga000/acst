.suckt  two_stage_single_output_op_amp_88_7 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mMainBias2 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mTelescopicFirstStageLoad3 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
mTelescopicFirstStageLoad4 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos
mTelescopicFirstStageLoad7 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mTelescopicFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos
mTelescopicFirstStageStageBias9 sourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos
mMainBias14 ibias ibias sourceNmos sourceNmos nmos
mMainBias15 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
mMainBias16 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_88_7

