** Name: two_stage_single_output_op_amp_101_3

.MACRO two_stage_single_output_op_amp_101_3 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=19e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=130e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=15e-6
mMainBias4 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=8e-6 W=326e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=19e-6
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=328e-6
mTelescopicFirstStageLoad8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=10e-6 W=38e-6
mMainBias9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=597e-6
mTelescopicFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=491e-6
mTelescopicFirstStageLoad11 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=8e-6 W=9e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=70e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=70e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=306e-6
mSecondStage1StageBias15 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=600e-6
mTelescopicFirstStageLoad16 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=8e-6 W=9e-6
mMainBias17 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=102e-6
mTelescopicFirstStageStageBias18 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=369e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.90001e-12
.EOM two_stage_single_output_op_amp_101_3

** Expected Performance Values: 
** Gain: 142 dB
** Power consumption: 4.65701 mW
** Area: 14942 (mu_m)^2
** Transit frequency: 2.55901 MHz
** Transit frequency with error factor: 2.55863 MHz
** Slew rate: 11.885 V/mu_s
** Phase margin: 60.1606°
** CMRR: 115 dB
** VoutMax: 4.03001 V
** VoutMin: 0.300001 V
** VcmMax: 3.21001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorNmos: 4.83334e+08 muA
** NormalTransistorPmos: -1.03414e+08 muA
** NormalTransistorPmos: -7.23899e+06 muA
** NormalTransistorPmos: -7.23899e+06 muA
** NormalTransistorNmos: 7.23801e+06 muA
** NormalTransistorNmos: 7.23801e+06 muA
** DiodeTransistorNmos: 7.23801e+06 muA
** NormalTransistorPmos: -4.97814e+08 muA
** NormalTransistorPmos: -4.97813e+08 muA
** NormalTransistorPmos: -7.23999e+06 muA
** NormalTransistorPmos: -7.23999e+06 muA
** NormalTransistorNmos: 3.10247e+08 muA
** NormalTransistorPmos: -3.10246e+08 muA
** NormalTransistorPmos: -3.10245e+08 muA
** DiodeTransistorNmos: 1.03415e+08 muA
** DiodeTransistorPmos: -4.83333e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.44101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.697001  V
** outVoltageBiasXXpXX1: 1.83401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21601  V
** innerSourceLoad2: 0.555001  V
** innerStageBias: 4.27901  V
** out1: 1.11001  V
** sourceGCC1: 2.99901  V
** sourceGCC2: 2.99601  V
** innerStageBias: 4.17501  V


.END