** Name: two_stage_single_output_op_amp_13_7

.MACRO two_stage_single_output_op_amp_13_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=11e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=7e-6 W=14e-6
mSimpleFirstStageTransconductor4 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=13e-6
mSimpleFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
mSecondStage1StageBias6 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=492e-6
mSimpleFirstStageTransconductor7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=13e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mSecondStage1Transconductor9 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=131e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=7e-6 W=14e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_13_7

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 2.37001 mW
** Area: 3481 (mu_m)^2
** Transit frequency: 2.50501 MHz
** Transit frequency with error factor: 2.50163 MHz
** Slew rate: 4.56442 V/mu_s
** Phase margin: 63.5984°
** CMRR: 93 dB
** negPSRR: 101 dB
** posPSRR: 88 dB
** VoutMax: 4.25 V
** VoutMin: 0.230001 V
** VcmMax: 3.54001 V
** VcmMin: 0.930001 V


** Expected Currents: 
** DiodeTransistorPmos: -1.02869e+07 muA
** NormalTransistorPmos: -1.02879e+07 muA
** NormalTransistorPmos: -1.02869e+07 muA
** DiodeTransistorPmos: -1.02879e+07 muA
** NormalTransistorNmos: 2.05731e+07 muA
** NormalTransistorNmos: 1.02861e+07 muA
** NormalTransistorNmos: 1.02861e+07 muA
** NormalTransistorNmos: 4.43365e+08 muA
** NormalTransistorPmos: -4.43364e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA


** Expected Voltages: 
** ibias: 0.636001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.23301  V
** innerTransistorStack1Load1: 4.23001  V
** out1: 3.13201  V
** sourceTransconductance: 1.80401  V


.END