** Name: symmetrical_op_amp192

.MACRO symmetrical_op_amp192 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=17e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=50e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=4e-6 W=10e-6
mSymmetricalFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=57e-6
mMainBias5 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=7e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=57e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=50e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
mSecondStage1StageBias10 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=6e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
mMainBias12 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=40e-6
mSymmetricalFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=23e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=23e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=54e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=9e-6 W=54e-6
mSymmetricalFirstStageLoad17 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=3e-6 W=122e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=3e-6 W=289e-6
mSecondStage1Transconductor19 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=289e-6
mSymmetricalFirstStageLoad20 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=122e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp192

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 0.722001 mW
** Area: 5121 (mu_m)^2
** Transit frequency: 2.78001 MHz
** Transit frequency with error factor: 2.78047 MHz
** Slew rate: 3.88671 V/mu_s
** Phase margin: 69.9009°
** CMRR: 135 dB
** negPSRR: 141 dB
** posPSRR: 62 dB
** VoutMax: 4.25 V
** VoutMin: 1.15001 V
** VcmMax: 4.81001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 2.35611e+07 muA
** NormalTransistorPmos: -1.64559e+07 muA
** NormalTransistorPmos: -1.64569e+07 muA
** NormalTransistorPmos: -1.64559e+07 muA
** NormalTransistorPmos: -1.64569e+07 muA
** NormalTransistorNmos: 3.29101e+07 muA
** DiodeTransistorNmos: 3.29111e+07 muA
** NormalTransistorNmos: 1.64551e+07 muA
** NormalTransistorNmos: 1.64551e+07 muA
** NormalTransistorNmos: 3.89891e+07 muA
** NormalTransistorNmos: 3.89881e+07 muA
** NormalTransistorPmos: -3.89899e+07 muA
** NormalTransistorPmos: -3.89889e+07 muA
** DiodeTransistorNmos: 3.89871e+07 muA
** DiodeTransistorNmos: 3.89861e+07 muA
** NormalTransistorPmos: -3.89879e+07 muA
** NormalTransistorPmos: -3.89889e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.35619e+07 muA


** Expected Voltages: 
** ibias: 1.14101  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 0.596001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 1.42901  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.571001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.87401  V
** innerStageBias: 0.468001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V
** inner: 0.569001  V


.END