.suckt  symmetrical_op_amp170 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m3 out2FirstStage out2FirstStage out1FirstStage out1FirstStage pmos
m4 out1FirstStage out1FirstStage sourcePmos sourcePmos pmos
m5 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage pmos
m6 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m7 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m8 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m9 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m10 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m11 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m12 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
m13 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m14 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m15 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
m16 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m18 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m19 ibias ibias sourceNmos sourceNmos nmos
m20 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end symmetrical_op_amp170

