.suckt  symmetrical_op_amp184 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 out2FirstStage ibias sourceNmos sourceNmos nmos
m3 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m4 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m5 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
m6 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m8 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m9 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m10 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m11 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m12 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m13 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
m14 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m16 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
m17 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m19 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m20 ibias ibias sourceNmos sourceNmos nmos
m21 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m22 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos
.end symmetrical_op_amp184

