.suckt  two_stage_single_output_op_amp_158_7 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m3 FirstStageYinnerLoad1 FirstStageYinnerLoad1 sourcePmos sourcePmos pmos
m4 outFirstStage FirstStageYinnerLoad1 sourcePmos sourcePmos pmos
m5 FirstStageYinnerLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m6 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m7 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m8 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m9 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m10 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m11 FirstStageYinnerLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c2 out sourceNmos 
m13 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m14 out outFirstStage sourcePmos sourcePmos pmos
m15 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m16 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m17 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_158_7

