** Name: two_stage_single_output_op_amp_147_8

.MACRO two_stage_single_output_op_amp_147_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=7e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=41e-6
mMainBias4 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=14e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=132e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=430e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=7e-6 W=541e-6
mSimpleFirstStageLoad11 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=7e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=132e-6
mSimpleFirstStageLoad13 FirstStageYinnerOutputLoad1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=184e-6
mMainBias14 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=405e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=359e-6
mSimpleFirstStageLoad16 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=184e-6
mMainBias17 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=229e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.2001e-12
.EOM two_stage_single_output_op_amp_147_8

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 11.3111 mW
** Area: 8315 (mu_m)^2
** Transit frequency: 6.48801 MHz
** Transit frequency with error factor: 6.47642 MHz
** Slew rate: 6.11495 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.25 V
** VoutMin: 0.75 V
** VcmMax: 5.25 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorPmos: -9.61939e+07 muA
** NormalTransistorPmos: -1.70884e+08 muA
** DiodeTransistorNmos: 4.49081e+07 muA
** DiodeTransistorNmos: 4.49091e+07 muA
** NormalTransistorNmos: 4.49081e+07 muA
** NormalTransistorNmos: 4.49091e+07 muA
** NormalTransistorPmos: -7.63359e+07 muA
** NormalTransistorPmos: -7.63359e+07 muA
** NormalTransistorNmos: 6.28531e+07 muA
** NormalTransistorNmos: 3.14271e+07 muA
** NormalTransistorNmos: 3.14271e+07 muA
** NormalTransistorNmos: 1.82254e+09 muA
** NormalTransistorNmos: 1.82254e+09 muA
** NormalTransistorPmos: -1.82253e+09 muA
** DiodeTransistorNmos: 9.61931e+07 muA
** DiodeTransistorNmos: 1.70885e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.628001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 1.15501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.13701  V
** innerTransistorStack2Load1: 1.13701  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.223001  V


.END