.suckt  symmetrical_op_amp76 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_FirstStage_Load_1 outFirstStage outFirstStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_StageBias_3 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_Symmetrical_FirstStage_StageBias_4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Transconductor_5 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_Symmetrical_FirstStage_Transconductor_6 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage2_StageBias_7 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos
m_Symmetrical_SecondStage2_StageBias_8 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage2_Transconductor_9 out outFirstStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_10 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_11 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_MainBias_12 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_Symmetrical_MainBias_13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
.end symmetrical_op_amp76

