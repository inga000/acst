** Name: one_stage_single_output_op_amp76

.MACRO one_stage_single_output_op_amp76 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=14e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=60e-6
m3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
m4 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=124e-6
m5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=24e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m7 out outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=12e-6
m8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=124e-6
m9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=19e-6
m10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=19e-6
m11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=60e-6
m12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=14e-6
m13 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=131e-6
m14 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
m15 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=412e-6
m16 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=131e-6
m17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=109e-6
m18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=109e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp76

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 3.36001 mW
** Area: 3515 (mu_m)^2
** Transit frequency: 2.73501 MHz
** Transit frequency with error factor: 2.73499 MHz
** Slew rate: 3.67786 V/mu_s
** Phase margin: 89.3815°
** CMRR: 143 dB
** VoutMax: 4.02001 V
** VoutMin: 0.430001 V
** VcmMax: 5.17001 V
** VcmMin: 1.78001 V


** Expected Currents: 
** NormalTransistorPmos: -1.71959e+07 muA
** NormalTransistorPmos: -4.13733e+08 muA
** NormalTransistorPmos: -7.36749e+07 muA
** NormalTransistorPmos: -1.1051e+08 muA
** NormalTransistorPmos: -7.36759e+07 muA
** NormalTransistorPmos: -1.10511e+08 muA
** DiodeTransistorNmos: 7.36741e+07 muA
** NormalTransistorNmos: 7.36751e+07 muA
** NormalTransistorNmos: 7.36741e+07 muA
** NormalTransistorNmos: 7.36731e+07 muA
** DiodeTransistorNmos: 7.36721e+07 muA
** NormalTransistorNmos: 3.68371e+07 muA
** NormalTransistorNmos: 3.68371e+07 muA
** DiodeTransistorNmos: 1.71951e+07 muA
** NormalTransistorNmos: 1.71941e+07 muA
** DiodeTransistorNmos: 4.13734e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.48201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outInputVoltageBiasXXnXX1: 1.56801  V
** outSourceVoltageBiasXXnXX1: 0.784001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 1.04001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.367001  V
** out1: 0.572001  V
** sourceGCC1: 4.22301  V
** sourceGCC2: 4.22301  V
** sourceTransconductance: 1.88001  V
** inner: 0.781001  V


.END