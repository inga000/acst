** Name: two_stage_single_output_op_amp_76_9

.MACRO two_stage_single_output_op_amp_76_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=55e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=420e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=319e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=46e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=422e-6
mMainBias6 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=5e-6 W=6e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=55e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=12e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=46e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=420e-6
mMainBias14 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=319e-6
mSecondStage1StageBias15 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=422e-6
mFoldedCascodeFirstStageLoad16 outFirstStage outVoltageBiasXXnXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=44e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=439e-6
mFoldedCascodeFirstStageLoad21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=24e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=255e-6
mMainBias23 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=548e-6
mMainBias24 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_76_9

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 8.39101 mW
** Area: 11633 (mu_m)^2
** Transit frequency: 4.24201 MHz
** Transit frequency with error factor: 4.24172 MHz
** Slew rate: 4.47576 V/mu_s
** Phase margin: 62.4525°
** CMRR: 138 dB
** VoutMax: 4.25 V
** VoutMin: 0.810001 V
** VcmMax: 5.17001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorPmos: -2.58538e+08 muA
** NormalTransistorPmos: -5.55604e+08 muA
** NormalTransistorPmos: -3.22929e+07 muA
** NormalTransistorPmos: -2.02109e+07 muA
** NormalTransistorPmos: -3.44709e+07 muA
** NormalTransistorPmos: -2.02109e+07 muA
** NormalTransistorPmos: -3.44709e+07 muA
** DiodeTransistorNmos: 2.02101e+07 muA
** NormalTransistorNmos: 2.02101e+07 muA
** NormalTransistorNmos: 2.02101e+07 muA
** NormalTransistorNmos: 2.85171e+07 muA
** DiodeTransistorNmos: 2.85161e+07 muA
** NormalTransistorNmos: 1.42591e+07 muA
** NormalTransistorNmos: 1.42591e+07 muA
** NormalTransistorNmos: 7.42891e+08 muA
** DiodeTransistorNmos: 7.4289e+08 muA
** NormalTransistorPmos: -7.4289e+08 muA
** DiodeTransistorNmos: 2.58539e+08 muA
** NormalTransistorNmos: 2.58538e+08 muA
** DiodeTransistorNmos: 5.55605e+08 muA
** NormalTransistorNmos: 5.55604e+08 muA
** DiodeTransistorNmos: 3.22921e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.15201  V
** outInputVoltageBiasXXnXX2: 1.21601  V
** outSourceVoltageBiasXXnXX1: 0.576001  V
** outSourceVoltageBiasXXnXX2: 0.608001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX3: 0.966001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.397001  V
** out1: 0.602001  V
** sourceGCC1: 4.17801  V
** sourceGCC2: 4.17801  V
** sourceTransconductance: 1.85701  V
** inner: 0.576001  V
** inner: 0.608001  V


.END