.suckt  two_stage_fully_differential_op_amp_51_12 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m3 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m4 outInputVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m5 outInputVoltageBiasXXnXX3 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m6 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m7 outFeedback outFeedback sourcePmos sourcePmos pmos
m8 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m9 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m14 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m15 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m16 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m17 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m18 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m19 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m20 out1 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m21 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m22 out1 outVoltageBiasXXpXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
m23 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m24 out2 outInputVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos
m25 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m26 out2 outVoltageBiasXXpXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
m27 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
m28 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m29 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m30 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
m31 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m32 outInputVoltageBiasXXnXX3 outInputVoltageBiasXXnXX3 VoltageBiasXXnXX3Yinner VoltageBiasXXnXX3Yinner nmos
m33 VoltageBiasXXnXX3Yinner outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m34 ibias ibias sourceNmos sourceNmos nmos
m35 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m36 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_51_12

