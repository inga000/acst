** Name: two_stage_single_output_op_amp_43_12

.MACRO two_stage_single_output_op_amp_43_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=16e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=5e-6 W=48e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=448e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=116e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=111e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=23e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=52e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=206e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=206e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=448e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=52e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=413e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=510e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=510e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=314e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=587e-6
mMainBias19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=121e-6
mMainBias20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=217e-6
mSecondStage1Transconductor21 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=594e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=111e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.8001e-12
.EOM two_stage_single_output_op_amp_43_12

** Expected Performance Values: 
** Gain: 136 dB
** Power consumption: 11.7901 mW
** Area: 14379 (mu_m)^2
** Transit frequency: 6.71801 MHz
** Transit frequency with error factor: 6.71237 MHz
** Slew rate: 5.51317 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** VoutMax: 4.25 V
** VoutMin: 0.800001 V
** VcmMax: 3.99001 V
** VcmMin: -0.339999 V


** Expected Currents: 
** NormalTransistorNmos: 3.45215e+08 muA
** NormalTransistorPmos: -5.25729e+07 muA
** NormalTransistorPmos: -9.58319e+07 muA
** NormalTransistorNmos: 1.03862e+08 muA
** NormalTransistorNmos: 1.73237e+08 muA
** NormalTransistorNmos: 1.03862e+08 muA
** NormalTransistorNmos: 1.73237e+08 muA
** DiodeTransistorPmos: -1.03861e+08 muA
** NormalTransistorPmos: -1.03861e+08 muA
** NormalTransistorPmos: -1.3875e+08 muA
** NormalTransistorPmos: -6.93759e+07 muA
** NormalTransistorPmos: -6.93759e+07 muA
** NormalTransistorNmos: 1.49797e+09 muA
** DiodeTransistorNmos: 1.49797e+09 muA
** NormalTransistorPmos: -1.49796e+09 muA
** NormalTransistorPmos: -1.49796e+09 muA
** DiodeTransistorNmos: 5.25721e+07 muA
** NormalTransistorNmos: 5.25731e+07 muA
** DiodeTransistorNmos: 9.58311e+07 muA
** DiodeTransistorNmos: 9.58301e+07 muA
** DiodeTransistorPmos: -3.45214e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.16501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.20601  V
** inputVoltageBiasXXnXX2: 1.37401  V
** out: 2.5  V
** outFirstStage: 4.06001  V
** outSourceVoltageBiasXXnXX1: 0.603001  V
** outSourceVoltageBiasXXnXX2: 0.627001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.03801  V
** sourceGCC1: 0.624001  V
** sourceGCC2: 0.624001  V
** sourceTransconductance: 3.23801  V
** innerTransconductance: 4.62401  V
** inner: 0.604001  V


.END