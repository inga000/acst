** Name: two_stage_single_output_op_amp_9_10

.MACRO two_stage_single_output_op_amp_9_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=317e-6
mSecondStage1StageBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=100e-6
mSimpleFirstStageTransconductor4 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=102e-6
mSimpleFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=55e-6
mSecondStage1StageBias6 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=550e-6
mSimpleFirstStageTransconductor7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=102e-6
mMainBias8 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=410e-6
mSimpleFirstStageLoad9 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=317e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=482e-6
mSecondStage1Transconductor11 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=4e-6 W=484e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.9001e-12
.EOM two_stage_single_output_op_amp_9_10

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 12.5871 mW
** Area: 9912 (mu_m)^2
** Transit frequency: 9.28001 MHz
** Transit frequency with error factor: 9.27397 MHz
** Slew rate: 10.3025 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** negPSRR: 107 dB
** posPSRR: 99 dB
** VoutMax: 4.25 V
** VoutMin: 0.340001 V
** VcmMax: 4.48001 V
** VcmMin: 0.920001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+09 muA
** NormalTransistorPmos: -6.73959e+07 muA
** NormalTransistorPmos: -6.73959e+07 muA
** DiodeTransistorPmos: -6.73959e+07 muA
** NormalTransistorNmos: 1.34792e+08 muA
** NormalTransistorNmos: 6.73951e+07 muA
** NormalTransistorNmos: 6.73951e+07 muA
** NormalTransistorNmos: 1.35721e+09 muA
** NormalTransistorPmos: -1.3572e+09 muA
** NormalTransistorPmos: -1.35721e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.01533e+09 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.04001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.24701  V
** out1: 3.50601  V
** sourceTransconductance: 1.91801  V
** innerTransconductance: 4.60401  V


.END