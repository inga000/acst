** Name: two_stage_single_output_op_amp_73_5

.MACRO two_stage_single_output_op_amp_73_5 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=119e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=26e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=5e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=7e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=396e-6
mMainBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=221e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=119e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=89e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=89e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=166e-6
mMainBias13 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=131e-6
mSecondStage1Transconductor14 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=219e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=6e-6 W=119e-6
mMainBias16 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=87e-6
mFoldedCascodeFirstStageLoad17 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=187e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mFoldedCascodeFirstStageLoad19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=7e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=396e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=187e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.70001e-12
.EOM two_stage_single_output_op_amp_73_5

** Expected Performance Values: 
** Gain: 133 dB
** Power consumption: 5.52801 mW
** Area: 14725 (mu_m)^2
** Transit frequency: 5.11701 MHz
** Transit frequency with error factor: 5.11734 MHz
** Slew rate: 4.29938 V/mu_s
** Phase margin: 60.1606°
** CMRR: 149 dB
** VoutMax: 3.17001 V
** VoutMin: 0.5 V
** VcmMax: 4.66001 V
** VcmMin: 1.28001 V


** Expected Currents: 
** NormalTransistorNmos: 1.65711e+07 muA
** NormalTransistorNmos: 2.50461e+07 muA
** NormalTransistorPmos: -3.77769e+07 muA
** NormalTransistorPmos: -5.89669e+07 muA
** NormalTransistorPmos: -3.77769e+07 muA
** NormalTransistorPmos: -5.89669e+07 muA
** NormalTransistorNmos: 3.77761e+07 muA
** NormalTransistorNmos: 3.77761e+07 muA
** DiodeTransistorNmos: 3.77761e+07 muA
** NormalTransistorNmos: 4.23771e+07 muA
** NormalTransistorNmos: 4.23761e+07 muA
** NormalTransistorNmos: 2.11891e+07 muA
** NormalTransistorNmos: 2.11891e+07 muA
** NormalTransistorNmos: 9.35992e+08 muA
** NormalTransistorPmos: -9.35991e+08 muA
** DiodeTransistorPmos: -9.35992e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.65719e+07 muA
** NormalTransistorPmos: -1.65729e+07 muA
** DiodeTransistorPmos: -2.50469e+07 muA
** DiodeTransistorPmos: -2.50459e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.37701  V
** out: 2.5  V
** outFirstStage: 0.905001  V
** outInputVoltageBiasXXpXX1: 2.60601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.80301  V
** outSourceVoltageBiasXXpXX2: 3.69101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerStageBias: 0.594001  V
** out1: 1.11001  V
** sourceGCC1: 3.09101  V
** sourceGCC2: 3.09101  V
** sourceTransconductance: 1.94501  V
** inner: 3.79801  V


.END