.suckt  two_stage_fully_differential_op_amp_38_1 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m3 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m5 outFeedback outFeedback sourceNmos sourceNmos nmos
m6 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m7 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
m8 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m9 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m14 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m15 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m16 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m17 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m18 out1FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m19 FirstStageYinnerTransistorStack1Load2 ibias sourcePmos sourcePmos pmos
m20 out2FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m21 FirstStageYinnerTransistorStack2Load2 ibias sourcePmos sourcePmos pmos
m22 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m23 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
m24 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m25 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m26 out1 out1FirstStage sourceNmos sourceNmos nmos
m27 out1 ibias sourcePmos sourcePmos pmos
m28 out2 out2FirstStage sourceNmos sourceNmos nmos
m29 out2 ibias sourcePmos sourcePmos pmos
m30 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m31 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m32 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m33 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_38_1

