** Name: two_stage_single_output_op_amp_195_9

.MACRO two_stage_single_output_op_amp_195_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=8e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=11e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=93e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=22e-6
m5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
m6 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=8e-6
m7 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=42e-6
m8 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=93e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=8e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=55e-6
m11 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=96e-6
m12 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
m13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=55e-6
m14 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=18e-6
m15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
m16 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=596e-6
m17 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=40e-6
m18 outFirstStage ibias sourcePmos sourcePmos pmos4 L=3e-6 W=290e-6
m19 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=589e-6
m20 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=290e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9e-12
.EOM two_stage_single_output_op_amp_195_9

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 7.59301 mW
** Area: 8595 (mu_m)^2
** Transit frequency: 4.89401 MHz
** Transit frequency with error factor: 4.88171 MHz
** Slew rate: 4.61234 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 1.19001 V
** VcmMax: 5.21001 V
** VcmMin: 1.59001 V


** Expected Currents: 
** NormalTransistorPmos: -1.40945e+08 muA
** NormalTransistorPmos: -9.60599e+06 muA
** DiodeTransistorNmos: 4.79791e+07 muA
** DiodeTransistorNmos: 4.79781e+07 muA
** NormalTransistorNmos: 4.79771e+07 muA
** NormalTransistorNmos: 4.79781e+07 muA
** NormalTransistorPmos: -6.89289e+07 muA
** NormalTransistorPmos: -6.89289e+07 muA
** NormalTransistorNmos: 4.19011e+07 muA
** NormalTransistorNmos: 4.19001e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** NormalTransistorNmos: 1.21029e+09 muA
** DiodeTransistorNmos: 1.21029e+09 muA
** NormalTransistorPmos: -1.21028e+09 muA
** DiodeTransistorNmos: 1.40946e+08 muA
** NormalTransistorNmos: 1.40947e+08 muA
** DiodeTransistorNmos: 9.60501e+06 muA
** DiodeTransistorNmos: 9.60401e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.23601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.31401  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.59201  V
** outSourceVoltageBiasXXnXX1: 0.796001  V
** outSourceVoltageBiasXXnXX2: 0.595001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.469001  V
** innerTransistorStack2Load1: 1.15601  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 0.797001  V


.END