.suckt  two_stage_single_output_op_amp_75_6 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_3 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_4 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_6 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m_SingleOutput_FirstStage_Load_7 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_8 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_9 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m_SingleOutput_FirstStage_Load_10 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_StageBias_11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_SingleOutput_FirstStage_StageBias_12 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Transconductor_13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_SingleOutput_FirstStage_Transconductor_14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_Transconductor_15 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_SingleOutput_SecondStage1_Transconductor_16 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_17 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_SingleOutput_SecondStage1_StageBias_18 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_19 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_20 ibias ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_21 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_SingleOutput_MainBias_22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_23 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m_SingleOutput_MainBias_24 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_75_6

