** Name: two_stage_single_output_op_amp_76_1

.MACRO two_stage_single_output_op_amp_76_1 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=121e-6
mMainBias2 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=15e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=48e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=253e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=25e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=190e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=121e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=105e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=105e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=253e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=15e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=468e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=168e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=192e-6
mMainBias15 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=482e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=574e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=120e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=120e-6
mMainBias19 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=148e-6
mSecondStage1StageBias20 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=536e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=574e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19e-12
.EOM two_stage_single_output_op_amp_76_1

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 9.99401 mW
** Area: 10962 (mu_m)^2
** Transit frequency: 8.23601 MHz
** Transit frequency with error factor: 8.23604 MHz
** Slew rate: 6.08044 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.69001 V
** VoutMin: 0.150001 V
** VcmMax: 5.10001 V
** VcmMin: 1.33001 V


** Expected Currents: 
** NormalTransistorNmos: 1.26917e+08 muA
** NormalTransistorNmos: 3.21133e+08 muA
** NormalTransistorPmos: -2.50145e+08 muA
** NormalTransistorPmos: -1.1656e+08 muA
** NormalTransistorPmos: -1.996e+08 muA
** NormalTransistorPmos: -1.1656e+08 muA
** NormalTransistorPmos: -1.996e+08 muA
** DiodeTransistorNmos: 1.16561e+08 muA
** NormalTransistorNmos: 1.16561e+08 muA
** NormalTransistorNmos: 1.16561e+08 muA
** NormalTransistorNmos: 1.66079e+08 muA
** DiodeTransistorNmos: 1.6608e+08 muA
** NormalTransistorNmos: 8.30391e+07 muA
** NormalTransistorNmos: 8.30391e+07 muA
** NormalTransistorNmos: 8.91366e+08 muA
** NormalTransistorPmos: -8.91365e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 2.50146e+08 muA
** DiodeTransistorPmos: -1.26916e+08 muA
** DiodeTransistorPmos: -3.21132e+08 muA


** Expected Voltages: 
** ibias: 1.16301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.958001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXnXX1: 0.582001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.13001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.351001  V
** out1: 0.556001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.92701  V
** inner: 0.580001  V


.END