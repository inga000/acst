** Name: two_stage_single_output_op_amp_190_9

.MACRO two_stage_single_output_op_amp_190_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=87e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=7e-6 W=84e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=30e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=407e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=25e-6
mSimpleFirstStageLoad9 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=30e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=87e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=84e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=407e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=8e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=25e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=103e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=103e-6
mSimpleFirstStageLoad18 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=52e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=328e-6
mSimpleFirstStageLoad20 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=52e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=45e-6
mMainBias22 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=137e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_190_9

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 5.38801 mW
** Area: 10522 (mu_m)^2
** Transit frequency: 3.22001 MHz
** Transit frequency with error factor: 3.21817 MHz
** Slew rate: 3.50001 V/mu_s
** Phase margin: 66.4632°
** CMRR: 118 dB
** VoutMax: 4.25 V
** VoutMin: 1.14001 V
** VcmMax: 4.84001 V
** VcmMin: 1.30001 V


** Expected Currents: 
** NormalTransistorPmos: -4.56239e+07 muA
** NormalTransistorPmos: -1.382e+08 muA
** NormalTransistorNmos: 9.59561e+07 muA
** NormalTransistorNmos: 9.59571e+07 muA
** DiodeTransistorNmos: 9.59561e+07 muA
** NormalTransistorPmos: -1.03871e+08 muA
** NormalTransistorPmos: -1.03872e+08 muA
** NormalTransistorPmos: -1.03872e+08 muA
** NormalTransistorPmos: -1.03872e+08 muA
** NormalTransistorNmos: 1.58301e+07 muA
** DiodeTransistorNmos: 1.58291e+07 muA
** NormalTransistorNmos: 7.91501e+06 muA
** NormalTransistorNmos: 7.91501e+06 muA
** NormalTransistorNmos: 6.66063e+08 muA
** DiodeTransistorNmos: 6.66062e+08 muA
** NormalTransistorPmos: -6.66062e+08 muA
** DiodeTransistorNmos: 4.56231e+07 muA
** NormalTransistorNmos: 4.56221e+07 muA
** DiodeTransistorNmos: 1.38201e+08 muA
** NormalTransistorNmos: 1.382e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.12601  V
** outInputVoltageBiasXXnXX2: 1.54401  V
** outSourceVoltageBiasXXnXX1: 0.563001  V
** outSourceVoltageBiasXXnXX2: 0.772001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.29501  V
** innerTransistorStack2Load1: 1.15501  V
** innerTransistorStack2Load2: 4.29501  V
** out1: 2.09501  V
** sourceTransconductance: 1.92201  V
** inner: 0.563001  V
** inner: 0.769001  V


.END