** Name: two_stage_single_output_op_amp_130_5

.MACRO two_stage_single_output_op_amp_130_5 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=13e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
m3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=4e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=558e-6
m5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=58e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=152e-6
m8 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=89e-6
m9 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=23e-6
m10 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=17e-6
m11 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=405e-6
m12 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=405e-6
m13 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=89e-6
m14 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=558e-6
m15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=7e-6 W=50e-6
m16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=29e-6
m17 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=8e-6 W=58e-6
m18 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=29e-6
m19 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=218e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.80001e-12
.EOM two_stage_single_output_op_amp_130_5

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 6.56801 mW
** Area: 12056 (mu_m)^2
** Transit frequency: 5.12801 MHz
** Transit frequency with error factor: 5.11717 MHz
** Slew rate: 24.2874 V/mu_s
** Phase margin: 60.1606°
** CMRR: 80 dB
** VoutMax: 3.32001 V
** VoutMin: 0.490001 V
** VcmMax: 3.51001 V
** VcmMin: -0.0899999 V


** Expected Currents: 
** NormalTransistorNmos: 7.34401e+06 muA
** NormalTransistorNmos: 5.46301e+06 muA
** NormalTransistorPmos: -7.25249e+07 muA
** NormalTransistorPmos: -7.25239e+07 muA
** DiodeTransistorPmos: -7.25249e+07 muA
** NormalTransistorNmos: 1.31414e+08 muA
** NormalTransistorNmos: 1.31413e+08 muA
** NormalTransistorNmos: 1.31413e+08 muA
** NormalTransistorNmos: 1.31413e+08 muA
** NormalTransistorPmos: -1.17778e+08 muA
** NormalTransistorPmos: -5.88889e+07 muA
** NormalTransistorPmos: -5.88889e+07 muA
** NormalTransistorNmos: 1.02792e+09 muA
** NormalTransistorPmos: -1.02791e+09 muA
** DiodeTransistorPmos: -1.02791e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.34499e+06 muA
** NormalTransistorPmos: -7.34599e+06 muA
** DiodeTransistorPmos: -5.46399e+06 muA


** Expected Voltages: 
** ibias: 1.19401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.897001  V
** outInputVoltageBiasXXpXX1: 2.75601  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outSourceVoltageBiasXXpXX1: 3.87801  V
** outVoltageBiasXXpXX2: 4.26201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.68601  V
** innerTransistorStack1Load2: 0.464001  V
** innerTransistorStack2Load2: 0.464001  V
** out1: 2.37201  V
** sourceTransconductance: 3.81401  V
** inner: 3.87301  V


.END