.suckt  two_stage_single_output_op_amp_85_1 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m3 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m4 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m5 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
m6 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos
m7 sourceTransconductance ibias sourcePmos sourcePmos pmos
m8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c2 out sourceNmos 
m10 out outFirstStage sourceNmos sourceNmos nmos
m11 out ibias sourcePmos sourcePmos pmos
m12 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m13 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
m14 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_85_1

