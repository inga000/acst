** Name: two_stage_single_output_op_amp_44_7

.MACRO two_stage_single_output_op_amp_44_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=39e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=431e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=92e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=149e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=149e-6
mSecondStage1StageBias8 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad9 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=92e-6
mFoldedCascodeFirstStageLoad10 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=431e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=49e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=49e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=455e-6
mMainBias14 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=156e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=461e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=290e-6
mMainBias17 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=433e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.40001e-12
.EOM two_stage_single_output_op_amp_44_7

** Expected Performance Values: 
** Gain: 110 dB
** Power consumption: 10.1291 mW
** Area: 9728 (mu_m)^2
** Transit frequency: 5.16301 MHz
** Transit frequency with error factor: 5.16311 MHz
** Slew rate: 18.4375 V/mu_s
** Phase margin: 60.1606°
** CMRR: 129 dB
** VoutMax: 4.25 V
** VoutMin: 0.150001 V
** VcmMax: 3.45001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.0953e+08 muA
** NormalTransistorPmos: -7.42819e+07 muA
** NormalTransistorNmos: 1.75227e+08 muA
** NormalTransistorNmos: 2.83791e+08 muA
** NormalTransistorNmos: 1.75227e+08 muA
** NormalTransistorNmos: 2.83791e+08 muA
** NormalTransistorPmos: -1.75226e+08 muA
** NormalTransistorPmos: -1.75226e+08 muA
** DiodeTransistorPmos: -1.75226e+08 muA
** NormalTransistorPmos: -2.1713e+08 muA
** NormalTransistorPmos: -1.08564e+08 muA
** NormalTransistorPmos: -1.08564e+08 muA
** NormalTransistorNmos: 1.15432e+09 muA
** NormalTransistorPmos: -1.15431e+09 muA
** DiodeTransistorNmos: 2.09531e+08 muA
** DiodeTransistorNmos: 7.42811e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.15201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 0.905001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.17401  V
** out1: 3.34901  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.76501  V


.END