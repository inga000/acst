** Name: two_stage_single_output_op_amp_170_3

.MACRO two_stage_single_output_op_amp_170_3 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=19e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=103e-6
m4 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=28e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=328e-6
m6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=41e-6
m7 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=7e-6 W=7e-6
m8 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=7e-6
m9 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=99e-6
m10 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=128e-6
m11 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=50e-6
m12 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=290e-6
m13 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=99e-6
m14 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=101e-6
m15 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=101e-6
m16 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=7e-6 W=7e-6
m17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=169e-6
m18 out outInputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=375e-6
m19 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=169e-6
m20 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=7e-6
m21 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=328e-6
m22 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=375e-6
m23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=103e-6
Capacitor1 outFirstStage out 17.9001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_170_3

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 7.54201 mW
** Area: 8158 (mu_m)^2
** Transit frequency: 3.00401 MHz
** Transit frequency with error factor: 3.00337 MHz
** Slew rate: 4.2427 V/mu_s
** Phase margin: 60.1606°
** CMRR: 77 dB
** VoutMax: 3.22001 V
** VoutMin: 0.340001 V
** VcmMax: 3.32001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 2.39121e+07 muA
** NormalTransistorNmos: 1.3814e+08 muA
** DiodeTransistorPmos: -9.95299e+06 muA
** DiodeTransistorPmos: -9.95399e+06 muA
** NormalTransistorPmos: -9.95299e+06 muA
** NormalTransistorPmos: -9.95399e+06 muA
** NormalTransistorNmos: 4.80911e+07 muA
** NormalTransistorNmos: 4.80921e+07 muA
** NormalTransistorNmos: 4.80911e+07 muA
** NormalTransistorNmos: 4.80921e+07 muA
** NormalTransistorPmos: -7.62789e+07 muA
** DiodeTransistorPmos: -7.62799e+07 muA
** NormalTransistorPmos: -3.81389e+07 muA
** NormalTransistorPmos: -3.81389e+07 muA
** NormalTransistorNmos: 1.24015e+09 muA
** NormalTransistorPmos: -1.24014e+09 muA
** NormalTransistorPmos: -1.24014e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.39129e+07 muA
** NormalTransistorPmos: -2.39139e+07 muA
** DiodeTransistorPmos: -1.38139e+08 muA
** DiodeTransistorPmos: -1.3814e+08 muA


** Expected Voltages: 
** ibias: 1.11701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.745001  V
** outInputVoltageBiasXXpXX1: 3.54801  V
** outInputVoltageBiasXXpXX2: 2.51501  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.27401  V
** outSourceVoltageBiasXXpXX2: 3.82501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.37201  V
** innerSourceLoad1: 3.68601  V
** innerTransistorStack1Load2: 0.560001  V
** innerTransistorStack2Load1: 3.67901  V
** innerTransistorStack2Load2: 0.560001  V
** sourceTransconductance: 3.28801  V
** innerStageBias: 3.68501  V
** inner: 4.27301  V


.END