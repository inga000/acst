** Name: one_stage_single_output_op_amp108

.MACRO one_stage_single_output_op_amp108 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=20e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mMainBias3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=37e-6
mTelescopicFirstStageStageBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=522e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=5e-6
mTelescopicFirstStageLoad6 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=69e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=69e-6
mTelescopicFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=69e-6
mTelescopicFirstStageLoad9 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=69e-6
mMainBias10 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mTelescopicFirstStageLoad11 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=61e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=452e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=452e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
mTelescopicFirstStageLoad15 out outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=61e-6
mMainBias16 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
mMainBias17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=240e-6
mTelescopicFirstStageStageBias18 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=522e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp108

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 1.20001 mW
** Area: 9562 (mu_m)^2
** Transit frequency: 6.70701 MHz
** Transit frequency with error factor: 6.70721 MHz
** Slew rate: 7.17366 V/mu_s
** Phase margin: 79.6412°
** CMRR: 147 dB
** VoutMax: 3.29001 V
** VoutMin: 0.300001 V
** VcmMax: 3.22001 V
** VcmMin: 0.0800001 V


** Expected Currents: 
** NormalTransistorNmos: 1.13451e+07 muA
** NormalTransistorPmos: -1.08089e+07 muA
** NormalTransistorPmos: -6.54119e+07 muA
** NormalTransistorPmos: -6.61829e+07 muA
** NormalTransistorPmos: -6.61849e+07 muA
** NormalTransistorNmos: 6.61821e+07 muA
** NormalTransistorNmos: 6.61831e+07 muA
** NormalTransistorNmos: 6.61841e+07 muA
** NormalTransistorNmos: 6.61831e+07 muA
** NormalTransistorPmos: -1.43712e+08 muA
** DiodeTransistorPmos: -1.43711e+08 muA
** NormalTransistorPmos: -6.61839e+07 muA
** NormalTransistorPmos: -6.61839e+07 muA
** DiodeTransistorNmos: 1.08081e+07 muA
** DiodeTransistorNmos: 6.54111e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.13459e+07 muA


** Expected Voltages: 
** ibias: 3.37601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.18901  V
** outVoltageBiasXXnXX0: 0.564001  V
** outVoltageBiasXXnXX1: 0.705001  V
** outVoltageBiasXXpXX2: 1.94501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.22001  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 3.00401  V
** sourceGCC2: 3.00401  V
** inner: 4.18501  V


.END