.suckt  two_stage_fully_differential_op_amp_19_3 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 outVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m5 outFeedback outFeedback sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m7 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m8 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m9 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m10 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m12 out1FirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m13 FirstStageYsourceGCC1 outFeedback sourcePmos sourcePmos pmos
m14 out2FirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m15 FirstStageYsourceGCC2 outFeedback sourcePmos sourcePmos pmos
m16 out1FirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m17 FirstStageYinnerTransistorStack1Load2 ibias sourceNmos sourceNmos nmos
m18 out2FirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m19 FirstStageYinnerTransistorStack2Load2 ibias sourceNmos sourceNmos nmos
m20 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m21 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m22 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m23 out1 out1FirstStage sourceNmos sourceNmos nmos
m24 out1 inputVoltageBiasXXpXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m25 SecondStage1YinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m26 out2 out2FirstStage sourceNmos sourceNmos nmos
m27 out2 inputVoltageBiasXXpXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m28 SecondStage2YinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m29 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m30 ibias ibias sourceNmos sourceNmos nmos
m31 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m32 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_19_3

