** Name: two_stage_single_output_op_amp_76_7

.MACRO two_stage_single_output_op_amp_76_7 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=19e-6
m2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=60e-6
m3 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
m4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=11e-6
m5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=51e-6
m6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=23e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=22e-6
m8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=19e-6
m9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=29e-6
m10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=29e-6
m11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=51e-6
m12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=11e-6
m13 out inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=395e-6
m14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=42e-6
m15 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=125e-6
m16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=55e-6
m17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=55e-6
m18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=487e-6
m19 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=58e-6
m20 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=504e-6
m21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=125e-6
m22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=8e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_76_7

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 6.74401 mW
** Area: 12206 (mu_m)^2
** Transit frequency: 3.36401 MHz
** Transit frequency with error factor: 3.36427 MHz
** Slew rate: 3.72146 V/mu_s
** Phase margin: 65.3172°
** CMRR: 143 dB
** VoutMax: 4.25 V
** VoutMin: 0.560001 V
** VcmMax: 5.13001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorPmos: -3.68499e+06 muA
** NormalTransistorPmos: -2.24394e+08 muA
** NormalTransistorPmos: -2.64329e+07 muA
** NormalTransistorPmos: -1.69219e+07 muA
** NormalTransistorPmos: -2.53909e+07 muA
** NormalTransistorPmos: -1.69219e+07 muA
** NormalTransistorPmos: -2.53909e+07 muA
** DiodeTransistorNmos: 1.69211e+07 muA
** NormalTransistorNmos: 1.69211e+07 muA
** NormalTransistorNmos: 1.69211e+07 muA
** NormalTransistorNmos: 1.69351e+07 muA
** DiodeTransistorNmos: 1.69341e+07 muA
** NormalTransistorNmos: 8.46801e+06 muA
** NormalTransistorNmos: 8.46801e+06 muA
** NormalTransistorNmos: 1.02347e+09 muA
** NormalTransistorPmos: -1.02346e+09 muA
** DiodeTransistorNmos: 3.68401e+06 muA
** NormalTransistorNmos: 3.68301e+06 muA
** DiodeTransistorNmos: 2.24395e+08 muA
** DiodeTransistorNmos: 2.64321e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.07301  V
** inputVoltageBiasXXnXX3: 0.961001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.16401  V
** outSourceVoltageBiasXXnXX1: 0.582001  V
** outSourceVoltageBiasXXpXX1: 4.15901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.655001  V
** innerTransistorStack2Load2: 0.450001  V
** sourceGCC1: 4.03801  V
** sourceGCC2: 4.03801  V
** sourceTransconductance: 1.91801  V
** inner: 0.581001  V


.END