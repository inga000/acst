.suckt  two_stage_fully_differential_op_amp_64_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_4 outVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_5 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_6 outFeedback outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m_FullyDifferential_FeedbackdStage_StageBias_8 FeedbackStageYinnerStageBias1 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m_FullyDifferential_FeedbackdStage_StageBias_10 FeedbackStageYinnerStageBias2 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackStage_Transconductor_11 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FeedbackStage_Transconductor_14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FirstStage_Load_15 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m_FullyDifferential_FirstStage_Load_16 FirstStageYsourceGCC1 outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_17 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m_FullyDifferential_FirstStage_Load_18 FirstStageYsourceGCC2 outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_19 out1FirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m_FullyDifferential_FirstStage_Load_20 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_21 out2FirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m_FullyDifferential_FirstStage_Load_22 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_StageBias_23 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_FullyDifferential_FirstStage_StageBias_24 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Transconductor_25 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_FullyDifferential_FirstStage_Transconductor_26 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_Transconductor_27 out1 inputVoltageBiasXXnXX2 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m_FullyDifferential_SecondStage1_Transconductor_28 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_29 out1 outVoltageBiasXXpXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m_FullyDifferential_SecondStage1_StageBias_30 SecondStage1YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_Transconductor_31 out2 inputVoltageBiasXXnXX2 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m_FullyDifferential_SecondStage2_Transconductor_32 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_StageBias_33 out2 outVoltageBiasXXpXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m_FullyDifferential_SecondStage2_StageBias_34 SecondStage2YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_35 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_FullyDifferential_MainBias_36 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_37 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_38 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_39 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_40 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_64_4

