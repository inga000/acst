.suckt  two_stage_fully_differential_op_amp_8_5 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 outVoltageBiasXXpXX3 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m4 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m5 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m6 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m7 outFeedback outFeedback sourceNmos sourceNmos nmos
m8 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX3 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m9 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
m10 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX3 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m11 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
m12 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m13 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m14 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m15 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m16 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m17 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m18 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m19 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m20 out1FirstStage outVoltageBiasXXpXX3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m21 FirstStageYinnerTransistorStack1Load2 ibias sourcePmos sourcePmos pmos
m22 out2FirstStage outVoltageBiasXXpXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m23 FirstStageYinnerTransistorStack2Load2 ibias sourcePmos sourcePmos pmos
m24 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m25 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m26 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m27 out1 out1FirstStage sourceNmos sourceNmos nmos
m28 out1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m29 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m30 out2 out2FirstStage sourceNmos sourceNmos nmos
m31 out2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m32 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m33 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m34 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m35 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m36 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m37 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m38 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m39 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m40 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_8_5

