** Name: two_stage_single_output_op_amp_61_10

.MACRO two_stage_single_output_op_amp_61_10 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=18e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=80e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=131e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=548e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=84e-6
m8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=177e-6
m9 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=84e-6
m10 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=108e-6
m11 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=108e-6
m12 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=511e-6
m13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=418e-6
m14 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=218e-6
m15 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=556e-6
m16 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=600e-6
m17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=131e-6
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=54e-6
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=54e-6
m20 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=410e-6
m21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=387e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 18.6001e-12
.EOM two_stage_single_output_op_amp_61_10

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 10.4061 mW
** Area: 10773 (mu_m)^2
** Transit frequency: 4.81001 MHz
** Transit frequency with error factor: 4.80993 MHz
** Slew rate: 6.58926 V/mu_s
** Phase margin: 60.1606°
** CMRR: 129 dB
** VoutMax: 4.27001 V
** VoutMin: 0.150001 V
** VcmMax: 3.18001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.40524e+08 muA
** NormalTransistorPmos: -1.13207e+08 muA
** NormalTransistorPmos: -1.52371e+08 muA
** NormalTransistorNmos: 1.23106e+08 muA
** NormalTransistorNmos: 2.05701e+08 muA
** NormalTransistorNmos: 1.23106e+08 muA
** NormalTransistorNmos: 2.05701e+08 muA
** DiodeTransistorPmos: -1.23105e+08 muA
** NormalTransistorPmos: -1.23105e+08 muA
** NormalTransistorPmos: -1.23105e+08 muA
** NormalTransistorPmos: -1.65186e+08 muA
** NormalTransistorPmos: -1.65185e+08 muA
** NormalTransistorPmos: -8.25939e+07 muA
** NormalTransistorPmos: -8.25939e+07 muA
** NormalTransistorNmos: 1.04374e+09 muA
** NormalTransistorPmos: -1.04373e+09 muA
** NormalTransistorPmos: -1.04373e+09 muA
** DiodeTransistorNmos: 1.13208e+08 muA
** DiodeTransistorNmos: 1.52372e+08 muA
** DiodeTransistorPmos: -3.40523e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.07601  V
** out: 2.5  V
** outFirstStage: 4.04601  V
** outVoltageBiasXXnXX2: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40001  V
** innerTransistorStack2Load2: 4.42701  V
** out1: 4.11101  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.35601  V
** innerTransconductance: 4.58701  V


.END