** Name: two_stage_single_output_op_amp_60_3

.MACRO two_stage_single_output_op_amp_60_3 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=13e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=83e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=8e-6 W=99e-6
m5 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=221e-6
m7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=20e-6
m9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=77e-6
m10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=77e-6
m11 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=198e-6
m12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=20e-6
m13 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
m14 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=74e-6
m15 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=83e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=124e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=124e-6
m18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=8e-6 W=221e-6
m19 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=261e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=99e-6
m21 out outInputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=121e-6
m22 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=9e-6 W=327e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_60_3

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 3.81601 mW
** Area: 14516 (mu_m)^2
** Transit frequency: 4.20701 MHz
** Transit frequency with error factor: 4.20712 MHz
** Slew rate: 4.26473 V/mu_s
** Phase margin: 63.0254°
** CMRR: 143 dB
** VoutMax: 3.51001 V
** VoutMin: 0.560001 V
** VcmMax: 3.31001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 8.76201e+06 muA
** NormalTransistorNmos: 2.82201e+07 muA
** NormalTransistorNmos: 1.94721e+07 muA
** NormalTransistorNmos: 2.93321e+07 muA
** NormalTransistorNmos: 1.94721e+07 muA
** NormalTransistorNmos: 2.93321e+07 muA
** NormalTransistorPmos: -1.94729e+07 muA
** NormalTransistorPmos: -1.94729e+07 muA
** DiodeTransistorPmos: -1.94729e+07 muA
** NormalTransistorPmos: -1.97229e+07 muA
** DiodeTransistorPmos: -1.97239e+07 muA
** NormalTransistorPmos: -9.86099e+06 muA
** NormalTransistorPmos: -9.86099e+06 muA
** NormalTransistorNmos: 6.57504e+08 muA
** NormalTransistorPmos: -6.57503e+08 muA
** NormalTransistorPmos: -6.57504e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -8.76299e+06 muA
** NormalTransistorPmos: -8.76399e+06 muA
** DiodeTransistorPmos: -2.82209e+07 muA
** DiodeTransistorPmos: -2.82199e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.968001  V
** outInputVoltageBiasXXpXX1: 3.47201  V
** outInputVoltageBiasXXpXX2: 3.09601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.23601  V
** outSourceVoltageBiasXXpXX2: 4.05901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.11101  V
** out1: 3.37301  V
** sourceGCC1: 0.527001  V
** sourceGCC2: 0.527001  V
** sourceTransconductance: 3.22701  V
** innerStageBias: 4.20901  V
** inner: 4.23501  V


.END