** Name: two_stage_single_output_op_amp_72_7

.MACRO two_stage_single_output_op_amp_72_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=63e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=40e-6
m3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=22e-6
m4 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
m5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=54e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=27e-6
m7 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=353e-6
m8 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
m9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
m10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
m11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=40e-6
m12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=63e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=400e-6
m14 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=5e-6 W=75e-6
m15 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=81e-6
m16 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=226e-6
m17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=5e-6 W=75e-6
m18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=74e-6
m19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=74e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_72_7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 7.72301 mW
** Area: 7691 (mu_m)^2
** Transit frequency: 3.71801 MHz
** Transit frequency with error factor: 3.71579 MHz
** Slew rate: 4.07698 V/mu_s
** Phase margin: 61.8795°
** CMRR: 98 dB
** VoutMax: 4.25 V
** VoutMin: 0.480001 V
** VcmMax: 5.08001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorPmos: -3.00479e+07 muA
** NormalTransistorPmos: -8.51199e+07 muA
** NormalTransistorPmos: -1.84439e+07 muA
** NormalTransistorPmos: -2.78709e+07 muA
** NormalTransistorPmos: -1.84439e+07 muA
** NormalTransistorPmos: -2.78709e+07 muA
** DiodeTransistorNmos: 1.84431e+07 muA
** NormalTransistorNmos: 1.84431e+07 muA
** NormalTransistorNmos: 1.88511e+07 muA
** DiodeTransistorNmos: 1.88501e+07 muA
** NormalTransistorNmos: 9.42601e+06 muA
** NormalTransistorNmos: 9.42601e+06 muA
** NormalTransistorNmos: 1.35379e+09 muA
** NormalTransistorPmos: -1.35378e+09 muA
** DiodeTransistorNmos: 3.00471e+07 muA
** NormalTransistorNmos: 3.00461e+07 muA
** DiodeTransistorNmos: 8.51191e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.14401  V
** outSourceVoltageBiasXXnXX1: 0.572001  V
** outSourceVoltageBiasXXpXX1: 4.11301  V
** outVoltageBiasXXnXX2: 0.881001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.870001  V
** sourceGCC1: 4.14701  V
** sourceGCC2: 4.14701  V
** sourceTransconductance: 1.91601  V
** inner: 0.571001  V


.END