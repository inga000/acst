** Name: symmetrical_op_amp42

.MACRO symmetrical_op_amp42 ibias in1 in2 out sourceNmos sourcePmos
m1 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=53e-6
m2 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=8e-6 W=91e-6
m3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=53e-6
m4 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=67e-6
m5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
m6 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=6e-6 W=67e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m8 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=8e-6 W=69e-6
m9 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=8e-6 W=69e-6
m10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=147e-6
m11 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=147e-6
m12 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=313e-6
m13 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=247e-6
m14 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=6e-6 W=67e-6
m15 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=313e-6
m16 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=67e-6
m17 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=34e-6
m18 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=67e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp42

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 2.63001 mW
** Area: 9390 (mu_m)^2
** Transit frequency: 7.26101 MHz
** Transit frequency with error factor: 7.26068 MHz
** Slew rate: 9.31818 V/mu_s
** Phase margin: 63.5984°
** CMRR: 141 dB
** negPSRR: 45 dB
** posPSRR: 48 dB
** VoutMax: 3.06001 V
** VoutMin: 0.510001 V
** VcmMax: 3.10001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorPmos: -2.50427e+08 muA
** DiodeTransistorNmos: 3.39641e+07 muA
** DiodeTransistorNmos: 3.39641e+07 muA
** NormalTransistorPmos: -6.79299e+07 muA
** NormalTransistorPmos: -6.79289e+07 muA
** NormalTransistorPmos: -3.39649e+07 muA
** NormalTransistorPmos: -3.39649e+07 muA
** NormalTransistorNmos: 9.33281e+07 muA
** NormalTransistorNmos: 9.33271e+07 muA
** NormalTransistorPmos: -9.33289e+07 muA
** DiodeTransistorPmos: -9.33299e+07 muA
** DiodeTransistorPmos: -9.42709e+07 muA
** NormalTransistorPmos: -9.42719e+07 muA
** NormalTransistorNmos: 9.42701e+07 muA
** NormalTransistorNmos: 9.42691e+07 muA
** DiodeTransistorNmos: 2.50428e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.913001  V
** inSourceStageBiasComplementarySecondStage: 3.74901  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 2.49801  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.29501  V
** sourceTransconductance: 3.27001  V
** innerTransconductance: 0.150001  V
** inner: 3.74601  V
** inner: 0.150001  V


.END