** Name: one_stage_single_output_op_amp60

.MACRO one_stage_single_output_op_amp60 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=54e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=105e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=84e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=584e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=52e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=75e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=75e-6
mFoldedCascodeFirstStageLoad9 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=52e-6
mFoldedCascodeFirstStageLoad10 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=105e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=84e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=84e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=584e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=84e-6
mMainBias15 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=455e-6
mFoldedCascodeFirstStageLoad16 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp60

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 1.42601 mW
** Area: 8456 (mu_m)^2
** Transit frequency: 3.66801 MHz
** Transit frequency with error factor: 3.66821 MHz
** Slew rate: 3.50001 V/mu_s
** Phase margin: 89.3815°
** CMRR: 130 dB
** VoutMax: 3.53001 V
** VoutMin: 0.770001 V
** VcmMax: 3.39001 V
** VcmMin: -0.379999 V


** Expected Currents: 
** NormalTransistorPmos: -5.41359e+07 muA
** NormalTransistorNmos: 7.00521e+07 muA
** NormalTransistorNmos: 1.05493e+08 muA
** NormalTransistorNmos: 7.00491e+07 muA
** NormalTransistorNmos: 1.0549e+08 muA
** NormalTransistorPmos: -7.00509e+07 muA
** NormalTransistorPmos: -7.00499e+07 muA
** DiodeTransistorPmos: -7.00509e+07 muA
** NormalTransistorPmos: -7.08819e+07 muA
** DiodeTransistorPmos: -7.08809e+07 muA
** NormalTransistorPmos: -3.54409e+07 muA
** NormalTransistorPmos: -3.54409e+07 muA
** DiodeTransistorNmos: 5.41351e+07 muA
** DiodeTransistorNmos: 5.41361e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.54301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.14601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.587001  V
** outSourceVoltageBiasXXpXX1: 4.27201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.16201  V
** out1: 2.96901  V
** sourceGCC1: 0.562001  V
** sourceGCC2: 0.562001  V
** sourceTransconductance: 3.21701  V
** inner: 4.27001  V


.END