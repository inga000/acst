** Name: two_stage_single_output_op_amp_60_9

.MACRO two_stage_single_output_op_amp_60_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=7e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=120e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=199e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=136e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=125e-6
mMainBias6 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=91e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=179e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=49e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=110e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=110e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mSecondStage1StageBias12 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=199e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=49e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=5e-6 W=125e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=33e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=33e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=179e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=91e-6
mMainBias19 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=225e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=333e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=72e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=8e-6 W=77e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.5e-12
.EOM two_stage_single_output_op_amp_60_9

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 4.29501 mW
** Area: 14736 (mu_m)^2
** Transit frequency: 3.12901 MHz
** Transit frequency with error factor: 3.129 MHz
** Slew rate: 3.59698 V/mu_s
** Phase margin: 60.1606°
** CMRR: 137 dB
** VoutMax: 4.25 V
** VoutMin: 1.32001 V
** VcmMax: 3.30001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.52129e+07 muA
** NormalTransistorPmos: -3.70049e+07 muA
** NormalTransistorNmos: 1.98991e+07 muA
** NormalTransistorNmos: 2.99301e+07 muA
** NormalTransistorNmos: 1.98991e+07 muA
** NormalTransistorNmos: 2.99301e+07 muA
** NormalTransistorPmos: -1.98999e+07 muA
** NormalTransistorPmos: -1.98999e+07 muA
** DiodeTransistorPmos: -1.98999e+07 muA
** NormalTransistorPmos: -2.00589e+07 muA
** DiodeTransistorPmos: -2.00579e+07 muA
** NormalTransistorPmos: -1.00299e+07 muA
** NormalTransistorPmos: -1.00299e+07 muA
** NormalTransistorNmos: 7.17022e+08 muA
** DiodeTransistorNmos: 7.17021e+08 muA
** NormalTransistorPmos: -7.17021e+08 muA
** DiodeTransistorNmos: 2.52121e+07 muA
** NormalTransistorNmos: 2.52111e+07 muA
** DiodeTransistorNmos: 3.70041e+07 muA
** DiodeTransistorNmos: 3.70051e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.48501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.73001  V
** inputVoltageBiasXXnXX2: 1.11901  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.865001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.24301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.22501  V
** out1: 3.32201  V
** sourceGCC1: 0.530001  V
** sourceGCC2: 0.530001  V
** sourceTransconductance: 3.24801  V
** inner: 0.862001  V
** inner: 4.24101  V


.END