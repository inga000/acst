.suckt  two_stage_fully_differential_op_amp_52_1 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 outInputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m3 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m4 outFeedback outFeedback sourcePmos sourcePmos pmos
m5 FeedbackStageYsourceTransconductance1 outInputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m6 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m7 FeedbackStageYsourceTransconductance2 outInputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m8 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m9 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m14 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m15 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m16 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m17 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m18 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m19 out1 out1FirstStage sourceNmos sourceNmos nmos
m20 out1 ibias sourcePmos sourcePmos pmos
m21 out2 out2FirstStage sourceNmos sourceNmos nmos
m22 out2 ibias sourcePmos sourcePmos pmos
m23 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m24 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m25 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m26 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m27 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_52_1

