** Name: two_stage_single_output_op_amp_38_7

.MACRO two_stage_single_output_op_amp_38_7 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=25e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=9e-6 W=15e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=32e-6
m4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
m5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=12e-6
m6 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=73e-6
m7 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=32e-6
m8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=15e-6
m9 out ibias sourceNmos sourceNmos nmos4 L=8e-6 W=600e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=73e-6
m11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=21e-6
m12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=71e-6
m13 FirstStageYinnerSourceLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=4e-6 W=214e-6
m14 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=57e-6
m15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=57e-6
m16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=555e-6
m17 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=214e-6
m18 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_38_7

** Expected Performance Values: 
** Gain: 103 dB
** Power consumption: 1.77701 mW
** Area: 10180 (mu_m)^2
** Transit frequency: 5.35201 MHz
** Transit frequency with error factor: 5.34865 MHz
** Slew rate: 5.04379 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** negPSRR: 163 dB
** posPSRR: 108 dB
** VoutMax: 4.84001 V
** VoutMin: 0.190001 V
** VcmMax: 5.14001 V
** VcmMin: 1.74001 V


** Expected Currents: 
** NormalTransistorNmos: 8.31601e+06 muA
** NormalTransistorNmos: 2.80711e+07 muA
** NormalTransistorPmos: -2.13569e+07 muA
** NormalTransistorPmos: -2.31739e+07 muA
** NormalTransistorPmos: -2.31749e+07 muA
** NormalTransistorPmos: -2.31739e+07 muA
** NormalTransistorPmos: -2.31749e+07 muA
** NormalTransistorNmos: 4.63451e+07 muA
** DiodeTransistorNmos: 4.63441e+07 muA
** NormalTransistorNmos: 2.31731e+07 muA
** NormalTransistorNmos: 2.31731e+07 muA
** NormalTransistorNmos: 2.41356e+08 muA
** NormalTransistorPmos: -2.41355e+08 muA
** DiodeTransistorNmos: 2.13561e+07 muA
** NormalTransistorNmos: 2.13561e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.31699e+06 muA
** DiodeTransistorPmos: -2.80719e+07 muA


** Expected Voltages: 
** ibias: 0.599001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.28001  V
** outInputVoltageBiasXXnXX1: 1.59201  V
** outSourceVoltageBiasXXnXX1: 0.796001  V
** outVoltageBiasXXpXX0: 4.27601  V
** outVoltageBiasXXpXX1: 3.71601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.17501  V
** innerTransistorStack1Load1: 4.43501  V
** innerTransistorStack2Load1: 4.43501  V
** sourceTransconductance: 1.94501  V
** inner: 0.796001  V


.END