** Name: one_stage_single_output_op_amp86

.MACRO one_stage_single_output_op_amp86 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=32e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=36e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=5e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=6e-6 W=32e-6
mTelescopicFirstStageLoad6 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=18e-6
mMainBias7 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=5e-6 W=267e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=172e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=172e-6
mTelescopicFirstStageLoad11 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=5e-6 W=267e-6
mMainBias12 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=10e-6
mTelescopicFirstStageStageBias13 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=271e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp86

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 0.496001 mW
** Area: 5149 (mu_m)^2
** Transit frequency: 3.77001 MHz
** Transit frequency with error factor: 3.77006 MHz
** Slew rate: 3.80583 V/mu_s
** Phase margin: 69.9009°
** CMRR: 153 dB
** VoutMax: 4.40001 V
** VoutMin: 0.840001 V
** VcmMax: 4.03001 V
** VcmMin: 0.480001 V


** Expected Currents: 
** NormalTransistorNmos: 2.80201e+06 muA
** NormalTransistorPmos: -2.81099e+06 muA
** NormalTransistorPmos: -3.68149e+07 muA
** NormalTransistorPmos: -3.68159e+07 muA
** NormalTransistorNmos: 3.68141e+07 muA
** NormalTransistorNmos: 3.68151e+07 muA
** DiodeTransistorNmos: 3.68141e+07 muA
** NormalTransistorPmos: -7.64319e+07 muA
** NormalTransistorPmos: -3.68149e+07 muA
** NormalTransistorPmos: -3.68149e+07 muA
** DiodeTransistorNmos: 2.81001e+06 muA
** DiodeTransistorPmos: -2.80299e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outVoltageBiasXXnXX0: 0.562001  V
** outVoltageBiasXXpXX1: 2.25801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21801  V
** innerTransistorStack2Load2: 0.690001  V
** out1: 1.25  V
** sourceGCC1: 3.01901  V
** sourceGCC2: 3.01901  V


.END