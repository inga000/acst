** Name: two_stage_single_output_op_amp_51_9

.MACRO two_stage_single_output_op_amp_51_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=28e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=554e-6
m3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=188e-6
m4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
m5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=35e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=25e-6
m7 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=554e-6
m8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=13e-6
m9 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=13e-6
m11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=13e-6
m12 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=10e-6 W=113e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=28e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=248e-6
m15 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=155e-6
m16 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=68e-6
m17 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=108e-6
m18 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=68e-6
m19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=97e-6
m20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=97e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.10001e-12
.EOM two_stage_single_output_op_amp_51_9

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 7.19401 mW
** Area: 12243 (mu_m)^2
** Transit frequency: 4.40801 MHz
** Transit frequency with error factor: 4.40763 MHz
** Slew rate: 4.21474 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 4.25 V
** VoutMin: 1.13001 V
** VcmMax: 5.11001 V
** VcmMin: 0.720001 V


** Expected Currents: 
** NormalTransistorPmos: -6.21139e+07 muA
** NormalTransistorPmos: -4.32789e+07 muA
** NormalTransistorPmos: -2.58059e+07 muA
** NormalTransistorPmos: -3.88709e+07 muA
** NormalTransistorPmos: -2.58059e+07 muA
** NormalTransistorPmos: -3.88709e+07 muA
** NormalTransistorNmos: 2.58051e+07 muA
** NormalTransistorNmos: 2.58051e+07 muA
** DiodeTransistorNmos: 2.58051e+07 muA
** NormalTransistorNmos: 2.61271e+07 muA
** NormalTransistorNmos: 1.30641e+07 muA
** NormalTransistorNmos: 1.30641e+07 muA
** NormalTransistorNmos: 1.23565e+09 muA
** DiodeTransistorNmos: 1.23565e+09 muA
** NormalTransistorPmos: -1.23564e+09 muA
** DiodeTransistorNmos: 6.21131e+07 muA
** NormalTransistorNmos: 6.21121e+07 muA
** DiodeTransistorNmos: 4.32781e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.53401  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.767001  V
** outSourceVoltageBiasXXpXX1: 4.13801  V
** outVoltageBiasXXnXX2: 0.570001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.706001  V
** out1: 1.26401  V
** sourceGCC1: 4.17601  V
** sourceGCC2: 4.17601  V
** sourceTransconductance: 1.94101  V
** inner: 0.766001  V


.END