** Name: two_stage_single_output_op_amp_203_8

.MACRO two_stage_single_output_op_amp_203_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=46e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=46e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=10e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=10e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=114e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=46e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=103e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=44e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mSecondStage1StageBias11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=116e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=46e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=103e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
mSimpleFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=418e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=516e-6
mSimpleFirstStageLoad17 outFirstStage outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=418e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.9001e-12
.EOM two_stage_single_output_op_amp_203_8

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 4.92801 mW
** Area: 10493 (mu_m)^2
** Transit frequency: 4.18701 MHz
** Transit frequency with error factor: 4.14217 MHz
** Slew rate: 3.94615 V/mu_s
** Phase margin: 60.1606°
** CMRR: 95 dB
** VoutMax: 4.84001 V
** VoutMin: 0.900001 V
** VcmMax: 5.02001 V
** VcmMin: 1.35001 V


** Expected Currents: 
** NormalTransistorNmos: 8.76201e+06 muA
** DiodeTransistorNmos: 3.46182e+08 muA
** NormalTransistorNmos: 3.46183e+08 muA
** NormalTransistorNmos: 3.46182e+08 muA
** DiodeTransistorNmos: 3.46183e+08 muA
** NormalTransistorPmos: -3.67979e+08 muA
** NormalTransistorPmos: -3.67979e+08 muA
** NormalTransistorNmos: 4.35951e+07 muA
** NormalTransistorNmos: 4.35941e+07 muA
** NormalTransistorNmos: 2.17981e+07 muA
** NormalTransistorNmos: 2.17981e+07 muA
** NormalTransistorNmos: 2.30865e+08 muA
** NormalTransistorNmos: 2.30864e+08 muA
** NormalTransistorPmos: -2.30864e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -8.76299e+06 muA


** Expected Voltages: 
** ibias: 1.20201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.27701  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 4.05101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.13901  V
** innerStageBias: 0.554001  V
** innerTransistorStack1Load1: 1.13901  V
** out1: 2.14301  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.453001  V


.END