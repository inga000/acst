.suckt  symmetrical_op_amp2 ibias in1 in2 out sourceNmos sourcePmos
m1 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos
m2 outFirstStage outFirstStage sourceNmos sourceNmos nmos
m3 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m4 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m5 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m6 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c1 out sourceNmos 
m7 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m9 out innerComplementarySecondStage sourcePmos sourcePmos pmos
m10 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos
m11 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m12 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m13 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m14 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp2

