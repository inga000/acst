** Name: symmetrical_op_amp80

.MACRO symmetrical_op_amp80 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=12e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=98e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=1e-6 W=65e-6
mSymmetricalFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mSecondStage1StageBias5 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad6 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=421e-6
mSymmetricalFirstStageLoad7 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=421e-6
mSymmetricalFirstStageStageBias8 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=600e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=98e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mMainBias11 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=120e-6
mSymmetricalFirstStageTransconductor12 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=115e-6
mSecondStage1StageBias13 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=107e-6
mSymmetricalFirstStageTransconductor14 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=115e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=535e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=535e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=600e-6
mSecondStage1Transconductor18 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp80

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 6.21801 mW
** Area: 7752 (mu_m)^2
** Transit frequency: 31.1301 MHz
** Transit frequency with error factor: 31.1304 MHz
** Slew rate: 31.7447 V/mu_s
** Phase margin: 61.8795°
** CMRR: 153 dB
** negPSRR: 81 dB
** posPSRR: 53 dB
** VoutMax: 4.65001 V
** VoutMin: 0.790001 V
** VcmMax: 4.66001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 9.97191e+07 muA
** DiodeTransistorPmos: -2.4711e+08 muA
** DiodeTransistorPmos: -2.4711e+08 muA
** NormalTransistorNmos: 4.9422e+08 muA
** DiodeTransistorNmos: 4.94219e+08 muA
** NormalTransistorNmos: 2.47111e+08 muA
** NormalTransistorNmos: 2.47111e+08 muA
** NormalTransistorNmos: 3.1988e+08 muA
** NormalTransistorNmos: 3.19879e+08 muA
** NormalTransistorPmos: -3.19879e+08 muA
** NormalTransistorPmos: -3.19878e+08 muA
** DiodeTransistorNmos: 3.19878e+08 muA
** DiodeTransistorNmos: 3.19877e+08 muA
** NormalTransistorPmos: -3.19877e+08 muA
** NormalTransistorPmos: -3.19878e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.97199e+07 muA


** Expected Voltages: 
** ibias: 1.15101  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceStageBiasComplementarySecondStage: 0.601001  V
** inSourceTransconductanceComplementarySecondStage: 4.25401  V
** innerComplementarySecondStage: 1.24601  V
** out: 2.5  V
** outFirstStage: 4.25401  V
** outSourceVoltageBiasXXnXX1: 0.576001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.93501  V
** innerStageBias: 0.653001  V
** innerTransconductance: 4.42201  V
** inner: 4.42201  V
** inner: 0.574001  V


.END