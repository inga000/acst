** Name: one_stage_single_output_op_amp97

.MACRO one_stage_single_output_op_amp97 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=46e-6
mTelescopicFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=70e-6
mTelescopicFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=70e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
mTelescopicFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=65e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=65e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=65e-6
mTelescopicFirstStageLoad9 out outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=65e-6
mMainBias10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mTelescopicFirstStageStageBias11 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=137e-6
mTelescopicFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=70e-6
mTelescopicFirstStageLoad13 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=70e-6
mMainBias14 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=152e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp97

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 0.840001 mW
** Area: 2287 (mu_m)^2
** Transit frequency: 3.27701 MHz
** Transit frequency with error factor: 3.27725 MHz
** Slew rate: 7.44594 V/mu_s
** Phase margin: 86.5167°
** CMRR: 149 dB
** VoutMax: 4.12001 V
** VoutMin: 0.530001 V
** VcmMax: 3.81001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorNmos: 8.77101e+06 muA
** NormalTransistorPmos: -8.73219e+07 muA
** NormalTransistorNmos: 3.09511e+07 muA
** NormalTransistorNmos: 3.09511e+07 muA
** DiodeTransistorPmos: -3.09519e+07 muA
** NormalTransistorPmos: -3.09529e+07 muA
** NormalTransistorPmos: -3.09519e+07 muA
** DiodeTransistorPmos: -3.09529e+07 muA
** NormalTransistorNmos: 1.49225e+08 muA
** NormalTransistorNmos: 3.09511e+07 muA
** NormalTransistorNmos: 3.09511e+07 muA
** DiodeTransistorNmos: 8.73211e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.77199e+06 muA


** Expected Voltages: 
** ibias: 0.633001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 4.25601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 4.27801  V
** innerTransistorStack1Load2: 4.27701  V
** out1: 3.55601  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END