** Name: two_stage_single_output_op_amp_162_1

.MACRO two_stage_single_output_op_amp_162_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=13e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=6e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=16e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=217e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=93e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=93e-6
mSimpleFirstStageLoad9 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=93e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=378e-6
mSimpleFirstStageLoad11 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=93e-6
mMainBias12 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=9e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=30e-6
mSimpleFirstStageTransconductor14 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=127e-6
mSimpleFirstStageLoad15 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=6e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=217e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=16e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=470e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=10e-6 W=12e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=127e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.90001e-12
.EOM two_stage_single_output_op_amp_162_1

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 4.31201 mW
** Area: 10014 (mu_m)^2
** Transit frequency: 2.88201 MHz
** Transit frequency with error factor: 2.88019 MHz
** Slew rate: 5.18301 V/mu_s
** Phase margin: 60.1606°
** CMRR: 81 dB
** VoutMax: 4.57001 V
** VoutMin: 0.380001 V
** VcmMax: 3.10001 V
** VcmMin: -0.259999 V


** Expected Currents: 
** NormalTransistorNmos: 3.42901e+06 muA
** NormalTransistorNmos: 1.15431e+07 muA
** NormalTransistorPmos: -1.21839e+07 muA
** NormalTransistorPmos: -1.21839e+07 muA
** DiodeTransistorPmos: -1.21839e+07 muA
** NormalTransistorNmos: 3.54271e+07 muA
** NormalTransistorNmos: 3.54271e+07 muA
** NormalTransistorNmos: 3.54271e+07 muA
** NormalTransistorNmos: 3.54271e+07 muA
** NormalTransistorPmos: -4.64889e+07 muA
** DiodeTransistorPmos: -4.64899e+07 muA
** NormalTransistorPmos: -2.32439e+07 muA
** NormalTransistorPmos: -2.32439e+07 muA
** NormalTransistorNmos: 7.66473e+08 muA
** NormalTransistorPmos: -7.66472e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.42999e+06 muA
** NormalTransistorPmos: -3.43099e+06 muA
** DiodeTransistorPmos: -1.15439e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.786001  V
** outInputVoltageBiasXXpXX1: 3.38001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19001  V
** outVoltageBiasXXpXX2: 4.00701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.68601  V
** innerTransistorStack1Load2: 0.618001  V
** innerTransistorStack2Load2: 0.618001  V
** out1: 2.37201  V
** sourceTransconductance: 3.34901  V
** inner: 4.18801  V


.END