** Name: symmetrical_op_amp51

.MACRO symmetrical_op_amp51 ibias in1 in2 out sourceNmos sourcePmos
m1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=73e-6
m3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
m4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=73e-6
m5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=10e-6
m6 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=92e-6
m8 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
m9 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=1e-6 W=22e-6
m10 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=1e-6 W=22e-6
m11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=164e-6
m12 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=164e-6
m13 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=126e-6
m14 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=326e-6
m15 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=3e-6 W=91e-6
m16 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m17 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=433e-6
m18 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=326e-6
m19 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=92e-6
m20 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=187e-6
m21 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=187e-6
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp51

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 2.36301 mW
** Area: 9766 (mu_m)^2
** Transit frequency: 6.55801 MHz
** Transit frequency with error factor: 6.55785 MHz
** Slew rate: 10.3625 V/mu_s
** Phase margin: 77.9223°
** CMRR: 148 dB
** negPSRR: 46 dB
** posPSRR: 54 dB
** VoutMax: 4.49001 V
** VoutMin: 0.390001 V
** VcmMax: 3.14001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 1.35361e+07 muA
** NormalTransistorPmos: -1.10269e+07 muA
** NormalTransistorPmos: -1.25562e+08 muA
** DiodeTransistorNmos: 4.66381e+07 muA
** DiodeTransistorNmos: 4.66381e+07 muA
** NormalTransistorPmos: -9.32769e+07 muA
** DiodeTransistorPmos: -9.32759e+07 muA
** NormalTransistorPmos: -4.66389e+07 muA
** NormalTransistorPmos: -4.66389e+07 muA
** NormalTransistorNmos: 1.04122e+08 muA
** NormalTransistorNmos: 1.04121e+08 muA
** NormalTransistorPmos: -1.04121e+08 muA
** NormalTransistorPmos: -1.04122e+08 muA
** NormalTransistorPmos: -1.05172e+08 muA
** NormalTransistorPmos: -1.05173e+08 muA
** NormalTransistorNmos: 1.05173e+08 muA
** NormalTransistorNmos: 1.05172e+08 muA
** DiodeTransistorNmos: 1.10261e+07 muA
** DiodeTransistorNmos: 1.25563e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.35369e+07 muA


** Expected Voltages: 
** ibias: 3.39601  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 3.68601  V
** inOutputTransconductanceComplementarySecondStage: 0.792001  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 4.12901  V
** inputVoltageBiasXXnXX0: 0.716001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.31601  V
** innerStageBias: 4.45001  V
** innerTransconductance: 0.150001  V
** inner: 4.68901  V
** inner: 0.150001  V
** inner: 4.19601  V


.END