** Name: two_stage_single_output_op_amp_46_8

.MACRO two_stage_single_output_op_amp_46_8 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=17e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=8e-6 W=153e-6
m4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=101e-6
m5 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=6e-6 W=106e-6
m6 out outInputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=125e-6
m7 outFirstStage outInputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
m8 FirstStageYout1 outInputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
m9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
m10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
m11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=171e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=82e-6
m13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=106e-6
m14 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=520e-6
m15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=101e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=37e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=37e-6
m18 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=8e-6 W=498e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_46_8

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 2.74501 mW
** Area: 12987 (mu_m)^2
** Transit frequency: 2.58701 MHz
** Transit frequency with error factor: 2.58705 MHz
** Slew rate: 5.07299 V/mu_s
** Phase margin: 61.3065°
** CMRR: 131 dB
** VoutMax: 4.25 V
** VoutMin: 0.770001 V
** VcmMax: 3.82001 V
** VcmMin: -0.389999 V


** Expected Currents: 
** NormalTransistorPmos: -3.39109e+07 muA
** NormalTransistorNmos: 2.29991e+07 muA
** NormalTransistorNmos: 3.94281e+07 muA
** NormalTransistorNmos: 2.29951e+07 muA
** NormalTransistorNmos: 3.94221e+07 muA
** DiodeTransistorPmos: -2.29979e+07 muA
** DiodeTransistorPmos: -2.29969e+07 muA
** NormalTransistorPmos: -2.29959e+07 muA
** NormalTransistorPmos: -2.29969e+07 muA
** NormalTransistorPmos: -3.28559e+07 muA
** NormalTransistorPmos: -1.64279e+07 muA
** NormalTransistorPmos: -1.64279e+07 muA
** NormalTransistorNmos: 4.16289e+08 muA
** NormalTransistorNmos: 4.16288e+08 muA
** NormalTransistorPmos: -4.16288e+08 muA
** DiodeTransistorNmos: 3.39101e+07 muA
** DiodeTransistorNmos: 3.39111e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.13301  V
** outSourceVoltageBiasXXnXX1: 0.575001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.15901  V
** innerTransistorStack2Load2: 4.15701  V
** out1: 3.32401  V
** sourceGCC1: 0.563001  V
** sourceGCC2: 0.563001  V
** sourceTransconductance: 3.50801  V
** innerStageBias: 0.529001  V


.END