** Name: one_stage_single_output_op_amp45

.MACRO one_stage_single_output_op_amp45 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=9e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
m3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=12e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=330e-6
m6 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
m7 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
m8 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=53e-6
m9 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=53e-6
m10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=175e-6
m11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=175e-6
m12 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=149e-6
m13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=330e-6
m14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=187e-6
m15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=187e-6
m16 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=137e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp45

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 1.29101 mW
** Area: 4807 (mu_m)^2
** Transit frequency: 4.01001 MHz
** Transit frequency with error factor: 4.0096 MHz
** Slew rate: 3.80665 V/mu_s
** Phase margin: 88.2356°
** CMRR: 144 dB
** VoutMax: 4.5 V
** VoutMin: 0.780001 V
** VcmMax: 3.93001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.26761e+07 muA
** NormalTransistorNmos: 6.67101e+06 muA
** NormalTransistorNmos: 7.62981e+07 muA
** NormalTransistorNmos: 1.14449e+08 muA
** NormalTransistorNmos: 7.62981e+07 muA
** NormalTransistorNmos: 1.14449e+08 muA
** DiodeTransistorPmos: -7.62989e+07 muA
** NormalTransistorPmos: -7.62989e+07 muA
** NormalTransistorPmos: -7.62989e+07 muA
** NormalTransistorPmos: -7.63029e+07 muA
** NormalTransistorPmos: -3.81509e+07 muA
** NormalTransistorPmos: -3.81509e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.26769e+07 muA
** DiodeTransistorPmos: -6.67199e+06 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** inputVoltageBiasXXpXX2: 4.08201  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.58701  V
** out1: 4.27501  V
** sourceGCC1: 0.529001  V
** sourceGCC2: 0.529001  V
** sourceTransconductance: 3.21501  V


.END