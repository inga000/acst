** Name: one_stage_single_output_op_amp73

.MACRO one_stage_single_output_op_amp73 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=8e-6
mMainBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=139e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=260e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=91e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=91e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=70e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=116e-6
mFoldedCascodeFirstStageLoad12 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=9e-6 W=30e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=301e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=374e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=374e-6
mFoldedCascodeFirstStageLoad16 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=301e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp73

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 2.52601 mW
** Area: 3564 (mu_m)^2
** Transit frequency: 9.15801 MHz
** Transit frequency with error factor: 9.158 MHz
** Slew rate: 6.08777 V/mu_s
** Phase margin: 86.5167°
** CMRR: 132 dB
** VoutMax: 4.11001 V
** VoutMin: 1.75 V
** VcmMax: 5.23001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorNmos: 7.73941e+07 muA
** NormalTransistorPmos: -1.22246e+08 muA
** NormalTransistorPmos: -2.08908e+08 muA
** NormalTransistorPmos: -1.22246e+08 muA
** NormalTransistorPmos: -2.08908e+08 muA
** NormalTransistorNmos: 1.22247e+08 muA
** NormalTransistorNmos: 1.22247e+08 muA
** DiodeTransistorNmos: 1.22247e+08 muA
** NormalTransistorNmos: 1.73322e+08 muA
** NormalTransistorNmos: 1.73321e+08 muA
** NormalTransistorNmos: 8.66611e+07 muA
** NormalTransistorNmos: 8.66611e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.73949e+07 muA
** DiodeTransistorPmos: -7.73959e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.25901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 1.09601  V
** innerStageBias: 0.471001  V
** out1: 2.15601  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.94501  V


.END