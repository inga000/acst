** Name: two_stage_single_output_op_amp_79_9

.MACRO two_stage_single_output_op_amp_79_9 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=9e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=315e-6
m3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=42e-6
m4 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=9e-6 W=18e-6
m5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=42e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=22e-6
m7 outFirstStage outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=42e-6
m8 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=315e-6
m9 FirstStageYinnerStageBias outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=9e-6 W=22e-6
m10 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=22e-6
m11 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=22e-6
m12 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=42e-6
m13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=7e-6
m14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=7e-6
m15 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=8e-6 W=79e-6
m16 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=9e-6
m17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=64e-6
m18 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=575e-6
m19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=51e-6
m20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=408e-6
m21 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=34e-6
m22 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=64e-6
m23 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=55e-6
m24 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=55e-6
Capacitor1 outFirstStage out 4.5e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_79_9

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 5.65201 mW
** Area: 14105 (mu_m)^2
** Transit frequency: 2.63301 MHz
** Transit frequency with error factor: 2.63253 MHz
** Slew rate: 3.52265 V/mu_s
** Phase margin: 67.0361°
** CMRR: 136 dB
** VoutMax: 4.25 V
** VoutMin: 1.34001 V
** VcmMax: 5.09001 V
** VcmMin: 1.51001 V


** Expected Currents: 
** NormalTransistorPmos: -2.35659e+07 muA
** NormalTransistorPmos: -1.86478e+08 muA
** NormalTransistorPmos: -1.54939e+07 muA
** NormalTransistorPmos: -1.59489e+07 muA
** NormalTransistorPmos: -2.54149e+07 muA
** NormalTransistorPmos: -1.59489e+07 muA
** NormalTransistorPmos: -2.54149e+07 muA
** NormalTransistorNmos: 1.59481e+07 muA
** NormalTransistorNmos: 1.59471e+07 muA
** NormalTransistorNmos: 1.59481e+07 muA
** NormalTransistorNmos: 1.59471e+07 muA
** NormalTransistorNmos: 1.89291e+07 muA
** NormalTransistorNmos: 1.89281e+07 muA
** NormalTransistorNmos: 9.46501e+06 muA
** NormalTransistorNmos: 9.46501e+06 muA
** NormalTransistorNmos: 8.34029e+08 muA
** DiodeTransistorNmos: 8.34028e+08 muA
** NormalTransistorPmos: -8.34028e+08 muA
** DiodeTransistorNmos: 2.35651e+07 muA
** NormalTransistorNmos: 2.35641e+07 muA
** DiodeTransistorNmos: 1.86479e+08 muA
** DiodeTransistorNmos: 1.54931e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.74201  V
** outSourceVoltageBiasXXnXX1: 0.871001  V
** outSourceVoltageBiasXXpXX1: 4.11601  V
** outVoltageBiasXXnXX2: 1.05601  V
** outVoltageBiasXXnXX3: 0.706001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.501001  V
** innerTransistorStack1Load2: 0.461001  V
** innerTransistorStack2Load2: 0.461001  V
** out1: 0.651001  V
** sourceGCC1: 4.12101  V
** sourceGCC2: 4.12101  V
** sourceTransconductance: 1.84101  V
** inner: 0.870001  V


.END