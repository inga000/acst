** Name: two_stage_single_output_op_amp_151_7

.MACRO two_stage_single_output_op_amp_151_7 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=18e-6
m2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=3e-6 W=6e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=11e-6
m5 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
m6 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
m7 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=6e-6
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=20e-6
m9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=20e-6
m11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=69e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=537e-6
m13 outFirstStage inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=83e-6
m14 FirstStageYout1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=83e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10.1001e-12
.EOM two_stage_single_output_op_amp_151_7

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 2.87501 mW
** Area: 5853 (mu_m)^2
** Transit frequency: 3.99101 MHz
** Transit frequency with error factor: 3.97396 MHz
** Slew rate: 3.76117 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.73001 V
** VoutMin: 0.180001 V
** VcmMax: 4.74001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorNmos: 1.44571e+07 muA
** DiodeTransistorNmos: 8.81081e+07 muA
** NormalTransistorNmos: 8.81081e+07 muA
** NormalTransistorNmos: 8.81081e+07 muA
** DiodeTransistorNmos: 8.81081e+07 muA
** NormalTransistorPmos: -1.07155e+08 muA
** NormalTransistorPmos: -1.07155e+08 muA
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 3.36148e+08 muA
** NormalTransistorPmos: -3.36147e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.44579e+07 muA


** Expected Voltages: 
** ibias: 0.586001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.77501  V
** out: 2.5  V
** outFirstStage: 4.17001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 1.13001  V
** innerTransistorStack2Load1: 1.13001  V
** out1: 2.26001  V
** sourceTransconductance: 1.94501  V


.END