** Name: two_stage_single_output_op_amp_30_12

.MACRO two_stage_single_output_op_amp_30_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=8e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=142e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=120e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=372e-6
mSimpleFirstStageLoad5 FirstStageYinnerLoad1 FirstStageYinnerLoad1 sourcePmos sourcePmos pmos4 L=10e-6 W=161e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=10e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=30e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=38e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=120e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=142e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=8e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
mSecondStage1StageBias13 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=372e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=38e-6
mMainBias15 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=62e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=553e-6
mSecondStage1Transconductor17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=4e-6 W=475e-6
mSimpleFirstStageLoad18 outFirstStage FirstStageYinnerLoad1 sourcePmos sourcePmos pmos4 L=10e-6 W=161e-6
mMainBias19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=26e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_30_12

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 3.03001 mW
** Area: 14957 (mu_m)^2
** Transit frequency: 5.62301 MHz
** Transit frequency with error factor: 5.61853 MHz
** Slew rate: 5.29953 V/mu_s
** Phase margin: 61.8795°
** CMRR: 100 dB
** negPSRR: 98 dB
** posPSRR: 91 dB
** VoutMax: 4.32001 V
** VoutMin: 0.890001 V
** VcmMax: 4.64001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 1.10561e+07 muA
** NormalTransistorNmos: 7.61491e+07 muA
** NormalTransistorPmos: -2.82269e+07 muA
** DiodeTransistorPmos: -1.20639e+07 muA
** NormalTransistorPmos: -1.20639e+07 muA
** NormalTransistorNmos: 2.41251e+07 muA
** DiodeTransistorNmos: 2.41241e+07 muA
** NormalTransistorNmos: 1.20631e+07 muA
** NormalTransistorNmos: 1.20631e+07 muA
** NormalTransistorNmos: 4.56478e+08 muA
** DiodeTransistorNmos: 4.56479e+08 muA
** NormalTransistorPmos: -4.56477e+08 muA
** NormalTransistorPmos: -4.56478e+08 muA
** DiodeTransistorNmos: 2.82261e+07 muA
** NormalTransistorNmos: 2.82261e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.10569e+07 muA
** DiodeTransistorPmos: -7.61499e+07 muA


** Expected Voltages: 
** ibias: 1.29201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.94101  V
** out: 2.5  V
** outFirstStage: 4.22101  V
** outInputVoltageBiasXXnXX1: 1.11801  V
** outSourceVoltageBiasXXnXX1: 0.559001  V
** outSourceVoltageBiasXXnXX2: 0.647001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad1: 4.23101  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.71201  V
** inner: 0.559001  V
** inner: 0.643001  V


.END