** Name: two_stage_single_output_op_amp_24_1

.MACRO two_stage_single_output_op_amp_24_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=28e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=253e-6
mSimpleFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=339e-6
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=8e-6 W=133e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=116e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=7e-6 W=116e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=291e-6
mSimpleFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=133e-6
mMainBias11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=28e-6
mSimpleFirstStageTransconductor12 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=181e-6
mSimpleFirstStageStageBias13 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=339e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=253e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=58e-6
mSecondStage1StageBias16 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=181e-6
mMainBias18 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=90e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_24_1

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 2.38501 mW
** Area: 13622 (mu_m)^2
** Transit frequency: 6.40301 MHz
** Transit frequency with error factor: 6.39757 MHz
** Slew rate: 6.89513 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** negPSRR: 107 dB
** posPSRR: 188 dB
** VoutMax: 4.84001 V
** VoutMin: 0.150001 V
** VcmMax: 3.20001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.79491e+07 muA
** NormalTransistorPmos: -4.15879e+07 muA
** NormalTransistorPmos: -2.68009e+07 muA
** NormalTransistorNmos: 3.16711e+07 muA
** NormalTransistorNmos: 3.16701e+07 muA
** NormalTransistorNmos: 3.16711e+07 muA
** NormalTransistorNmos: 3.16701e+07 muA
** NormalTransistorPmos: -6.33449e+07 muA
** DiodeTransistorPmos: -6.33459e+07 muA
** NormalTransistorPmos: -3.16719e+07 muA
** NormalTransistorPmos: -3.16719e+07 muA
** NormalTransistorNmos: 2.77249e+08 muA
** NormalTransistorPmos: -2.77248e+08 muA
** DiodeTransistorNmos: 4.15871e+07 muA
** DiodeTransistorNmos: 2.68001e+07 muA
** DiodeTransistorPmos: -4.79499e+07 muA
** NormalTransistorPmos: -4.79509e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.37001  V
** outSourceVoltageBiasXXpXX1: 4.18501  V
** outVoltageBiasXXnXX0: 0.607001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.23501  V
** inner: 4.18501  V


.END