.suckt  two_stage_fully_differential_op_amp_50_7 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_3 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_4 outFeedback outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_5 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX1 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m_FullyDifferential_FeedbackdStage_StageBias_6 FeedbackStageYinnerStageBias1 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX1 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m_FullyDifferential_FeedbackdStage_StageBias_8 FeedbackStageYinnerStageBias2 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackStage_Transconductor_9 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_11 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FeedbackStage_Transconductor_12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FirstStage_Load_13 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_14 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_StageBias_15 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_FullyDifferential_FirstStage_StageBias_16 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Transconductor_17 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_FullyDifferential_FirstStage_Transconductor_18 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_StageBias_19 out1 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_Transconductor_20 out1 out1FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_StageBias_21 out2 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_Transconductor_22 out2 out2FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_23 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_24 ibias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_25 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_50_7

