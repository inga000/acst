** Name: one_stage_single_output_op_amp51

.MACRO one_stage_single_output_op_amp51 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=76e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=16e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=72e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=76e-6
mFoldedCascodeFirstStageTransconductor6 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=138e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=138e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=182e-6
mMainBias9 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=75e-6
mFoldedCascodeFirstStageLoad10 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=98e-6
mFoldedCascodeFirstStageLoad11 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=475e-6
mFoldedCascodeFirstStageLoad12 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=238e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=238e-6
mFoldedCascodeFirstStageLoad14 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=475e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp51

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 3.56401 mW
** Area: 4829 (mu_m)^2
** Transit frequency: 10.4391 MHz
** Transit frequency with error factor: 10.4387 MHz
** Slew rate: 9.57873 V/mu_s
** Phase margin: 86.5167°
** CMRR: 147 dB
** VoutMax: 4.02001 V
** VoutMin: 1.01001 V
** VcmMax: 5.14001 V
** VcmMin: 0.850001 V


** Expected Currents: 
** NormalTransistorNmos: 9.28471e+07 muA
** NormalTransistorPmos: -1.92913e+08 muA
** NormalTransistorPmos: -3.04939e+08 muA
** NormalTransistorPmos: -1.92913e+08 muA
** NormalTransistorPmos: -3.04939e+08 muA
** NormalTransistorNmos: 1.92914e+08 muA
** NormalTransistorNmos: 1.92914e+08 muA
** DiodeTransistorNmos: 1.92914e+08 muA
** NormalTransistorNmos: 2.24052e+08 muA
** NormalTransistorNmos: 1.12026e+08 muA
** NormalTransistorNmos: 1.12026e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.28479e+07 muA
** DiodeTransistorPmos: -9.28489e+07 muA


** Expected Voltages: 
** ibias: 0.676001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.16701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.861001  V
** out1: 1.41801  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.92501  V


.END