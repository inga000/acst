** Name: two_stage_single_output_op_amp_31_8

.MACRO two_stage_single_output_op_amp_31_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=5e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
mSimpleFirstStageStageBias4 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=19e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=465e-6
mSecondStage1StageBias8 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=228e-6
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=19e-6
mSimpleFirstStageLoad10 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
mSecondStage1Transconductor11 out outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=229e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=4e-6 W=37e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_31_8

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 2.46301 mW
** Area: 3099 (mu_m)^2
** Transit frequency: 2.91701 MHz
** Transit frequency with error factor: 2.91398 MHz
** Slew rate: 3.592 V/mu_s
** Phase margin: 60.1606°
** CMRR: 104 dB
** negPSRR: 97 dB
** posPSRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 0.780001 V
** VcmMax: 4.37001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorPmos: -8.82999e+06 muA
** NormalTransistorPmos: -8.82999e+06 muA
** DiodeTransistorPmos: -8.82999e+06 muA
** NormalTransistorNmos: 1.76571e+07 muA
** NormalTransistorNmos: 1.76581e+07 muA
** NormalTransistorNmos: 8.82901e+06 muA
** NormalTransistorNmos: 8.82901e+06 muA
** NormalTransistorNmos: 4.65026e+08 muA
** NormalTransistorNmos: 4.65025e+08 muA
** NormalTransistorPmos: -4.65025e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA


** Expected Voltages: 
** ibias: 1.18001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.19401  V
** innerStageBias: 0.570001  V
** out1: 3.39801  V
** sourceTransconductance: 1.89801  V
** innerStageBias: 0.555001  V


.END