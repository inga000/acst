** Name: two_stage_single_output_op_amp_37_8

.MACRO two_stage_single_output_op_amp_37_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=10e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
m3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m4 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=102e-6
m5 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=241e-6
m6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=20e-6
m7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=22e-6
m8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=20e-6
m9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=23e-6
m10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=464e-6
m11 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=151e-6
m12 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=27e-6
m13 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=7e-6 W=12e-6
m14 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=7e-6 W=12e-6
m15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=27e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_37_8

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 2.97701 mW
** Area: 2789 (mu_m)^2
** Transit frequency: 3.13201 MHz
** Transit frequency with error factor: 3.12894 MHz
** Slew rate: 4.74889 V/mu_s
** Phase margin: 60.1606°
** CMRR: 94 dB
** negPSRR: 94 dB
** posPSRR: 90 dB
** VoutMax: 4.29001 V
** VoutMin: 0.770001 V
** VcmMax: 4.81001 V
** VcmMin: 1.35001 V


** Expected Currents: 
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -1.09529e+07 muA
** NormalTransistorPmos: -1.09539e+07 muA
** NormalTransistorPmos: -1.09529e+07 muA
** NormalTransistorPmos: -1.09539e+07 muA
** NormalTransistorNmos: 2.19041e+07 muA
** NormalTransistorNmos: 2.19031e+07 muA
** NormalTransistorNmos: 1.09521e+07 muA
** NormalTransistorNmos: 1.09521e+07 muA
** NormalTransistorNmos: 4.61874e+08 muA
** NormalTransistorNmos: 4.61873e+08 muA
** NormalTransistorPmos: -4.61873e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.72301  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.561001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** out1: 3.83601  V
** sourceTransconductance: 1.85301  V
** innerStageBias: 0.498001  V


.END