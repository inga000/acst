** Name: one_stage_single_output_op_amp93

.MACRO one_stage_single_output_op_amp93 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=6e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=15e-6
mTelescopicFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
mTelescopicFirstStageLoad5 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=44e-6
mTelescopicFirstStageTransconductor6 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=74e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=74e-6
mTelescopicFirstStageLoad8 out outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=44e-6
mMainBias9 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=6e-6
mTelescopicFirstStageStageBias10 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=57e-6
mTelescopicFirstStageLoad11 FirstStageYout1 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mTelescopicFirstStageLoad12 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=62e-6
mMainBias13 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=19e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp93

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 0.571001 mW
** Area: 1511 (mu_m)^2
** Transit frequency: 2.98601 MHz
** Transit frequency with error factor: 2.98624 MHz
** Slew rate: 4.69729 V/mu_s
** Phase margin: 88.2356°
** CMRR: 152 dB
** VoutMax: 3.94001 V
** VoutMin: 0.580001 V
** VcmMax: 4.19001 V
** VcmMin: 0.830001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00551e+07 muA
** NormalTransistorPmos: -3.77169e+07 muA
** NormalTransistorNmos: 2.81891e+07 muA
** NormalTransistorNmos: 2.81881e+07 muA
** NormalTransistorPmos: -2.81899e+07 muA
** NormalTransistorPmos: -2.81889e+07 muA
** DiodeTransistorPmos: -2.81899e+07 muA
** NormalTransistorNmos: 9.40931e+07 muA
** NormalTransistorNmos: 2.81891e+07 muA
** NormalTransistorNmos: 2.81891e+07 muA
** DiodeTransistorNmos: 3.77161e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.00559e+07 muA


** Expected Voltages: 
** ibias: 0.685001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 3.76701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 4.09901  V
** out1: 3.375  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END