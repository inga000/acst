** Name: two_stage_single_output_op_amp_34_9

.MACRO two_stage_single_output_op_amp_34_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=7e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=24e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=17e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=525e-6
mSimpleFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=13e-6
mMainBias6 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=21e-6
mMainBias7 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=379e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=22e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=17e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=24e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mMainBias12 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mSecondStage1StageBias13 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=525e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=22e-6
mMainBias15 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=303e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=13e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=114e-6
mSimpleFirstStageLoad18 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=5e-6 W=129e-6
mMainBias19 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=26e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_34_9

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 6.32501 mW
** Area: 8261 (mu_m)^2
** Transit frequency: 4.89401 MHz
** Transit frequency with error factor: 4.89086 MHz
** Slew rate: 4.61201 V/mu_s
** Phase margin: 65.3172°
** CMRR: 98 dB
** negPSRR: 155 dB
** posPSRR: 96 dB
** VoutMax: 4.40001 V
** VoutMin: 0.770001 V
** VcmMax: 4.09001 V
** VcmMin: 1.60001 V


** Expected Currents: 
** NormalTransistorNmos: 4.25228e+08 muA
** NormalTransistorNmos: 4.26431e+07 muA
** NormalTransistorPmos: -2.93319e+07 muA
** DiodeTransistorPmos: -1.04769e+07 muA
** NormalTransistorPmos: -1.04769e+07 muA
** NormalTransistorPmos: -1.04769e+07 muA
** NormalTransistorNmos: 2.09511e+07 muA
** DiodeTransistorNmos: 2.09501e+07 muA
** NormalTransistorNmos: 1.04761e+07 muA
** NormalTransistorNmos: 1.04761e+07 muA
** NormalTransistorNmos: 7.36779e+08 muA
** DiodeTransistorNmos: 7.3678e+08 muA
** NormalTransistorPmos: -7.36778e+08 muA
** DiodeTransistorNmos: 2.93311e+07 muA
** NormalTransistorNmos: 2.93301e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -4.25227e+08 muA
** DiodeTransistorPmos: -4.26439e+07 muA


** Expected Voltages: 
** ibias: 1.17501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.83601  V
** outInputVoltageBiasXXnXX1: 1.44601  V
** outSourceVoltageBiasXXnXX1: 0.723001  V
** outSourceVoltageBiasXXnXX2: 0.588001  V
** outVoltageBiasXXpXX0: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.40001  V
** out1: 3.83601  V
** sourceTransconductance: 1.94501  V
** inner: 0.722001  V
** inner: 0.586001  V


.END