.suckt  symmetrical_op_amp122 ibias in1 in2 out sourceNmos sourcePmos
m1 out1FirstStage out1FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m2 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
m3 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m4 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m6 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m7 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m8 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m9 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m10 out out1FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m11 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m12 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos
m13 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m14 innerComplementarySecondStage inSourceTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m15 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m16 ibias ibias sourceNmos sourceNmos nmos
.end symmetrical_op_amp122

