** Name: two_stage_single_output_op_amp_29_9

.MACRO two_stage_single_output_op_amp_29_9 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=5e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=22e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=230e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
m6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=111e-6
m7 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=230e-6
m8 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=30e-6
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=46e-6
m10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
m11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=46e-6
m12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=217e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=22e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=566e-6
m15 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=111e-6
m16 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=49e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.60001e-12
.EOM two_stage_single_output_op_amp_29_9

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 5.67001 mW
** Area: 5822 (mu_m)^2
** Transit frequency: 11.3641 MHz
** Transit frequency with error factor: 11.3008 MHz
** Slew rate: 28.033 V/mu_s
** Phase margin: 60.1606°
** CMRR: 86 dB
** negPSRR: 126 dB
** posPSRR: 84 dB
** VoutMax: 4.73001 V
** VoutMin: 0.800001 V
** VcmMax: 4.57001 V
** VcmMin: 1.82001 V


** Expected Currents: 
** NormalTransistorNmos: 1.42851e+07 muA
** NormalTransistorPmos: -7.08339e+07 muA
** DiodeTransistorPmos: -1.4429e+08 muA
** NormalTransistorPmos: -1.4429e+08 muA
** NormalTransistorNmos: 2.8858e+08 muA
** NormalTransistorNmos: 2.88579e+08 muA
** NormalTransistorNmos: 1.44291e+08 muA
** NormalTransistorNmos: 1.44291e+08 muA
** NormalTransistorNmos: 7.50316e+08 muA
** DiodeTransistorNmos: 7.50315e+08 muA
** NormalTransistorPmos: -7.50315e+08 muA
** DiodeTransistorNmos: 7.08331e+07 muA
** NormalTransistorNmos: 7.08341e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.42859e+07 muA


** Expected Voltages: 
** ibias: 1.26601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.03501  V
** out: 2.5  V
** outFirstStage: 4.16501  V
** outInputVoltageBiasXXnXX1: 1.20201  V
** outSourceVoltageBiasXXnXX1: 0.601001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.610001  V
** out1: 4.16501  V
** sourceTransconductance: 1.48401  V
** inner: 0.602001  V


.END