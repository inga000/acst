.suckt  two_stage_single_output_op_amp_14_8 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m_SingleOutput_FirstStage_Load_4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerOutputLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_5 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_SingleOutput_FirstStage_Load_6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerOutputLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_StageBias_7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Transconductor_8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_SingleOutput_FirstStage_Transconductor_9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_StageBias_10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m_SingleOutput_SecondStage1_StageBias_11 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_Transconductor_12 out outFirstStage sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_13 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_14 ibias ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_15 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_14_8

