.suckt  two_stage_single_output_op_amp_138_9 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mMainBias2 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mSimpleFirstStageLoad3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad5 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad7 FirstStageYinnerOutputLoad1 inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor12 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias14 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
mSecondStage1StageBias15 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos
mMainBias17 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
mMainBias18 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias19 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
mMainBias20 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias21 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_138_9

