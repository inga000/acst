** Name: symmetrical_op_amp50

.MACRO symmetrical_op_amp50 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=39e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=25e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=2e-6 W=10e-6
mSymmetricalFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=144e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=32e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=32e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=2e-6 W=19e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=19e-6
mSymmetricalFirstStageStageBias12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=144e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=25e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=39e-6
mMainBias15 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=160e-6
mSymmetricalFirstStageTransconductor16 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=81e-6
mSecondStage1StageBias17 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=210e-6
mSymmetricalFirstStageTransconductor18 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=81e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp50

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 0.980001 mW
** Area: 3230 (mu_m)^2
** Transit frequency: 4.92501 MHz
** Transit frequency with error factor: 4.92471 MHz
** Slew rate: 4.87756 V/mu_s
** Phase margin: 85.3708°
** CMRR: 150 dB
** negPSRR: 52 dB
** posPSRR: 64 dB
** VoutMax: 3.81001 V
** VoutMin: 0.440001 V
** VcmMax: 3.23001 V
** VcmMin: 0.0300001 V


** Expected Currents: 
** NormalTransistorPmos: -4.08229e+07 muA
** DiodeTransistorNmos: 1.87141e+07 muA
** DiodeTransistorNmos: 1.87141e+07 muA
** NormalTransistorPmos: -3.74299e+07 muA
** DiodeTransistorPmos: -3.74289e+07 muA
** NormalTransistorPmos: -1.87149e+07 muA
** NormalTransistorPmos: -1.87149e+07 muA
** NormalTransistorNmos: 4.89201e+07 muA
** NormalTransistorNmos: 4.89211e+07 muA
** NormalTransistorPmos: -4.89209e+07 muA
** NormalTransistorPmos: -4.89219e+07 muA
** DiodeTransistorPmos: -4.89229e+07 muA
** DiodeTransistorPmos: -4.89239e+07 muA
** NormalTransistorNmos: 4.89221e+07 muA
** NormalTransistorNmos: 4.89211e+07 muA
** DiodeTransistorNmos: 4.08221e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.842001  V
** inSourceStageBiasComplementarySecondStage: 3.96601  V
** inSourceTransconductanceComplementarySecondStage: 0.596001  V
** innerComplementarySecondStage: 2.65901  V
** out: 2.5  V
** outFirstStage: 0.596001  V
** outSourceVoltageBiasXXpXX1: 4.19601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.22501  V
** innerStageBias: 3.38401  V
** innerTransconductance: 0.191001  V
** inner: 0.191001  V
** inner: 4.19301  V


.END