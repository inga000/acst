.suckt  two_stage_fully_differential_op_amp_66_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m2 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m5 outFeedback outFeedback sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance1 outVoltageBiasXXnXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m7 FeedbackStageYinnerStageBias1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m8 FeedbackStageYsourceTransconductance2 outVoltageBiasXXnXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m9 FeedbackStageYinnerStageBias2 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m14 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m15 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m16 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m17 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m18 sourceTransconductance outVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m19 FirstStageYinnerStageBias inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m20 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m21 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m22 out1 outVoltageBiasXXnXX2 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m23 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m24 out1 ibias SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m25 SecondStage1YinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m26 out2 outVoltageBiasXXnXX2 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m27 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m28 out2 ibias SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m29 SecondStage2YinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m30 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
m31 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m32 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m33 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m34 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_66_4

