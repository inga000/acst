.suckt  two_stage_fully_differential_op_amp_59_2 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 outVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
m5 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m6 outFeedback outFeedback sourcePmos sourcePmos pmos
m7 FeedbackStageYsourceTransconductance1 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m8 FeedbackStageYsourceTransconductance2 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m9 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m14 FirstStageYsourceGCC1 outFeedback sourcePmos sourcePmos pmos
m15 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m16 FirstStageYsourceGCC2 outFeedback sourcePmos sourcePmos pmos
m17 out1FirstStage outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m18 out2FirstStage outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m19 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m20 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m21 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m22 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m23 out1 outVoltageBiasXXnXX2 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m24 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m25 out1 ibias sourcePmos sourcePmos pmos
m26 out2 outVoltageBiasXXnXX2 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m27 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m28 out2 ibias sourcePmos sourcePmos pmos
m29 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m30 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m31 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m32 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m33 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m34 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_59_2

