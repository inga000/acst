.suckt  two_stage_single_output_op_amp_129_4 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m5 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos
m6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m7 FirstStageYout1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m8 outFirstStage outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m9 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c2 out sourceNmos 
m12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m13 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m14 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m15 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos
m16 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m17 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m18 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m19 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_129_4

