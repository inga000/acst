** Name: two_stage_single_output_op_amp_114_10

.MACRO two_stage_single_output_op_amp_114_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=19e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=306e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=95e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=177e-6
mSecondStage1StageBias7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=23e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=23e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=23e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=6e-6 W=501e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=23e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=256e-6
mMainBias15 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=6e-6 W=600e-6
mTelescopicFirstStageStageBias16 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=306e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=346e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=599e-6
mTelescopicFirstStageLoad19 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mMainBias20 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=17e-6
mMainBias21 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=242e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.80001e-12
.EOM two_stage_single_output_op_amp_114_10

** Expected Performance Values: 
** Gain: 104 dB
** Power consumption: 5.99401 mW
** Area: 14348 (mu_m)^2
** Transit frequency: 5.33401 MHz
** Transit frequency with error factor: 5.32997 MHz
** Slew rate: 12.6473 V/mu_s
** Phase margin: 60.1606°
** CMRR: 86 dB
** VoutMax: 4.59001 V
** VoutMin: 0.220001 V
** VcmMax: 4.47001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 1.71791e+08 muA
** NormalTransistorNmos: 4.02635e+08 muA
** NormalTransistorPmos: -1.67759e+07 muA
** NormalTransistorPmos: -2.38864e+08 muA
** NormalTransistorNmos: 1.46031e+07 muA
** NormalTransistorNmos: 1.46031e+07 muA
** DiodeTransistorPmos: -1.46039e+07 muA
** NormalTransistorPmos: -1.46039e+07 muA
** NormalTransistorNmos: 2.6807e+08 muA
** DiodeTransistorNmos: 2.68069e+08 muA
** NormalTransistorNmos: 1.46031e+07 muA
** NormalTransistorNmos: 1.46031e+07 muA
** NormalTransistorNmos: 3.29544e+08 muA
** NormalTransistorPmos: -3.29543e+08 muA
** NormalTransistorPmos: -3.29544e+08 muA
** DiodeTransistorNmos: 1.67751e+07 muA
** NormalTransistorNmos: 1.67741e+07 muA
** DiodeTransistorNmos: 2.38865e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.7179e+08 muA
** DiodeTransistorPmos: -4.02634e+08 muA


** Expected Voltages: 
** ibias: 0.622001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.20401  V
** outInputVoltageBiasXXnXX1: 1.16201  V
** outSourceVoltageBiasXXnXX1: 0.581001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 3.86301  V
** outVoltageBiasXXpXX1: 2.92801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.21601  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 3.66701  V
** inner: 0.580001  V


.END