** Name: two_stage_single_output_op_amp_5_5

.MACRO two_stage_single_output_op_amp_5_5 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=18e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=10e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=42e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=10e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=520e-6
m6 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=554e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=271e-6
m8 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=46e-6
m9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=101e-6
m10 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=101e-6
m11 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=8e-6 W=271e-6
m12 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=71e-6
m13 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=520e-6
m14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=141e-6
m15 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=19e-6
m16 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=141e-6
m17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=536e-6
m18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_5_5

** Expected Performance Values: 
** Gain: 108 dB
** Power consumption: 6.23301 mW
** Area: 10046 (mu_m)^2
** Transit frequency: 27.6971 MHz
** Transit frequency with error factor: 27.6777 MHz
** Slew rate: 27.8508 V/mu_s
** Phase margin: 65.3172°
** CMRR: 106 dB
** negPSRR: 108 dB
** posPSRR: 233 dB
** VoutMax: 3.76001 V
** VoutMin: 0.150001 V
** VcmMax: 4.05001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.06201e+07 muA
** NormalTransistorPmos: -4.54999e+06 muA
** NormalTransistorPmos: -1.69939e+07 muA
** NormalTransistorNmos: 6.45331e+07 muA
** NormalTransistorNmos: 6.45341e+07 muA
** NormalTransistorNmos: 6.45351e+07 muA
** NormalTransistorNmos: 6.45341e+07 muA
** NormalTransistorPmos: -1.29066e+08 muA
** NormalTransistorPmos: -6.45339e+07 muA
** NormalTransistorPmos: -6.45339e+07 muA
** NormalTransistorNmos: 1.05538e+09 muA
** NormalTransistorPmos: -1.05537e+09 muA
** DiodeTransistorPmos: -1.05537e+09 muA
** DiodeTransistorNmos: 4.54901e+06 muA
** DiodeTransistorNmos: 1.69931e+07 muA
** DiodeTransistorPmos: -2.06209e+07 muA
** NormalTransistorPmos: -2.06209e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.20501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.19601  V
** outSourceVoltageBiasXXpXX1: 4.09801  V
** outVoltageBiasXXnXX0: 0.598001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.22401  V
** inner: 4.09801  V


.END