** Name: two_stage_single_output_op_amp_4_4

.MACRO two_stage_single_output_op_amp_4_4 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=35e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=36e-6
mSecondStage1StageBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=25e-6
mMainBias4 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=62e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=28e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=56e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=36e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=10e-6 W=238e-6
mSecondStage1Transconductor9 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=87e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=35e-6
mMainBias11 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=506e-6
mSimpleFirstStageTransconductor12 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=15e-6
mSimpleFirstStage_StageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=151e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=597e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=545e-6
mSecondStage1StageBias16 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=540e-6
mSimpleFirstStageTransconductor17 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=15e-6
mMainBias18 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=193e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_4_4

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 5.60901 mW
** Area: 14824 (mu_m)^2
** Transit frequency: 2.70401 MHz
** Transit frequency with error factor: 2.69479 MHz
** Slew rate: 8.81796 V/mu_s
** Phase margin: 61.3065°
** CMRR: 92 dB
** negPSRR: 86 dB
** posPSRR: 88 dB
** VoutMax: 4.57001 V
** VoutMin: 0.75 V
** VcmMax: 3.44001 V
** VcmMin: 0.580001 V


** Expected Currents: 
** NormalTransistorNmos: 5.63381e+08 muA
** NormalTransistorPmos: -7.02459e+07 muA
** NormalTransistorPmos: -1.95911e+08 muA
** DiodeTransistorNmos: 2.74791e+07 muA
** DiodeTransistorNmos: 2.74781e+07 muA
** NormalTransistorNmos: 2.74791e+07 muA
** NormalTransistorNmos: 2.74781e+07 muA
** NormalTransistorPmos: -5.49589e+07 muA
** NormalTransistorPmos: -2.74799e+07 muA
** NormalTransistorPmos: -2.74799e+07 muA
** NormalTransistorNmos: 2.17228e+08 muA
** NormalTransistorNmos: 2.17227e+08 muA
** NormalTransistorPmos: -2.17227e+08 muA
** NormalTransistorPmos: -2.17228e+08 muA
** DiodeTransistorNmos: 7.02451e+07 muA
** DiodeTransistorNmos: 1.95912e+08 muA
** DiodeTransistorPmos: -5.6338e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.15201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.15401  V
** out: 2.5  V
** outFirstStage: 0.735001  V
** outVoltageBiasXXnXX0: 0.731001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 1.14001  V
** innerSourceLoad1: 0.569001  V
** innerTransistorStack2Load1: 0.568001  V
** sourceTransconductance: 3.77701  V
** innerStageBias: 4.40001  V
** innerTransconductance: 0.330001  V


.END