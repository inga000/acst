** Name: two_stage_single_output_op_amp_60_5

.MACRO two_stage_single_output_op_amp_60_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=13e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=141e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=17e-6
mMainBias5 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=4e-6 W=15e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=63e-6
mSecondStage1StageBias7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=528e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=20e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=77e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=77e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=87e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=20e-6
mMainBias13 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=14e-6
mMainBias14 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=87e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=141e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=61e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=61e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=63e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=17e-6
mMainBias20 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=15e-6
mSecondStage1StageBias21 out outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=4e-6 W=528e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=7e-6 W=65e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_60_5

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 6.31401 mW
** Area: 9097 (mu_m)^2
** Transit frequency: 4.21601 MHz
** Transit frequency with error factor: 4.21619 MHz
** Slew rate: 4.3088 V/mu_s
** Phase margin: 72.7657°
** CMRR: 136 dB
** VoutMax: 3.03001 V
** VoutMin: 0.560001 V
** VcmMax: 3.06001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 5.33301e+06 muA
** NormalTransistorNmos: 3.31411e+07 muA
** NormalTransistorNmos: 1.94721e+07 muA
** NormalTransistorNmos: 2.93321e+07 muA
** NormalTransistorNmos: 1.94721e+07 muA
** NormalTransistorNmos: 2.93321e+07 muA
** NormalTransistorPmos: -1.94729e+07 muA
** NormalTransistorPmos: -1.94729e+07 muA
** DiodeTransistorPmos: -1.94729e+07 muA
** NormalTransistorPmos: -1.97229e+07 muA
** DiodeTransistorPmos: -1.97239e+07 muA
** NormalTransistorPmos: -9.86099e+06 muA
** NormalTransistorPmos: -9.86099e+06 muA
** NormalTransistorNmos: 1.15562e+09 muA
** NormalTransistorPmos: -1.15561e+09 muA
** DiodeTransistorPmos: -1.15561e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.33399e+06 muA
** NormalTransistorPmos: -5.33499e+06 muA
** DiodeTransistorPmos: -3.31419e+07 muA
** NormalTransistorPmos: -3.31429e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.968001  V
** outInputVoltageBiasXXpXX1: 3.22201  V
** outInputVoltageBiasXXpXX2: 2.46601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.11101  V
** outSourceVoltageBiasXXpXX2: 3.73301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.26001  V
** out1: 3.35201  V
** sourceGCC1: 0.527001  V
** sourceGCC2: 0.527001  V
** sourceTransconductance: 3.22801  V
** inner: 4.10901  V
** inner: 3.73001  V


.END