** Name: two_stage_single_output_op_amp_197_9

.MACRO two_stage_single_output_op_amp_197_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=33e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=44e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=30e-6
mMainBias4 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=8e-6 W=29e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=416e-6
mMainBias6 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=119e-6
mMainBias7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=64e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=33e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=38e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=8e-6 W=25e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=30e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=416e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=44e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=38e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=400e-6
mSimpleFirstStageLoad18 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=400e-6
mSimpleFirstStageLoad19 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=600e-6
mMainBias20 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
mMainBias21 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=38e-6
mSecondStage1Transconductor22 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=529e-6
mSimpleFirstStageLoad23 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=600e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_197_9

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 9.07001 mW
** Area: 9233 (mu_m)^2
** Transit frequency: 4.67001 MHz
** Transit frequency with error factor: 4.66634 MHz
** Slew rate: 4.40127 V/mu_s
** Phase margin: 63.0254°
** CMRR: 126 dB
** VoutMax: 4.25 V
** VoutMin: 0.720001 V
** VcmMax: 4.98001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorPmos: -6.45979e+07 muA
** NormalTransistorPmos: -3.77649e+07 muA
** DiodeTransistorNmos: 3.87904e+08 muA
** DiodeTransistorNmos: 3.87905e+08 muA
** NormalTransistorNmos: 3.87904e+08 muA
** NormalTransistorNmos: 3.87905e+08 muA
** NormalTransistorPmos: -3.98243e+08 muA
** NormalTransistorPmos: -3.98244e+08 muA
** NormalTransistorPmos: -3.98243e+08 muA
** NormalTransistorPmos: -3.98244e+08 muA
** NormalTransistorNmos: 2.06791e+07 muA
** NormalTransistorNmos: 2.06781e+07 muA
** NormalTransistorNmos: 1.03401e+07 muA
** NormalTransistorNmos: 1.03401e+07 muA
** NormalTransistorNmos: 8.95192e+08 muA
** DiodeTransistorNmos: 8.95191e+08 muA
** NormalTransistorPmos: -8.95191e+08 muA
** DiodeTransistorNmos: 6.45971e+07 muA
** NormalTransistorNmos: 6.45961e+07 muA
** DiodeTransistorNmos: 3.77641e+07 muA
** DiodeTransistorNmos: 3.77631e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.12801  V
** inputVoltageBiasXXnXX2: 1.33401  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.564001  V
** outSourceVoltageBiasXXnXX2: 0.579001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15401  V
** innerStageBias: 0.649001  V
** innerTransistorStack1Load2: 4.15401  V
** innerTransistorStack2Load1: 1.15401  V
** innerTransistorStack2Load2: 4.15401  V
** out1: 2.20701  V
** sourceTransconductance: 1.94501  V
** inner: 0.563001  V


.END