.suckt  two_stage_single_output_op_amp_130_2 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mMainBias2 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad4 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad8 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1Transconductor13 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mSecondStage1Transconductor14 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias15 out ibias sourcePmos sourcePmos pmos
mMainBias16 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias17 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias18 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_130_2

