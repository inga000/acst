** Name: symmetrical_op_amp67

.MACRO symmetrical_op_amp67 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=13e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=159e-6
mSymmetricalFirstStageLoad5 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=159e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=7e-6
mSymmetricalFirstStageStageBias7 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=534e-6
mSymmetricalFirstStageStageBias8 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=118e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=39e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias10 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=39e-6
mMainBias11 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos4 L=5e-6 W=133e-6
mSymmetricalFirstStageTransconductor12 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=52e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias13 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=1e-6 W=74e-6
mSecondStage1StageBias14 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=73e-6
mSymmetricalFirstStageTransconductor15 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=52e-6
mMainBias16 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=15e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=148e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=148e-6
mMainBias19 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=90e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor20 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=475e-6
mSecondStage1Transconductor21 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=475e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp67

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 5.33401 mW
** Area: 9175 (mu_m)^2
** Transit frequency: 4.96601 MHz
** Transit frequency with error factor: 4.96617 MHz
** Slew rate: 19.1224 V/mu_s
** Phase margin: 72.1927°
** CMRR: 132 dB
** negPSRR: 45 dB
** posPSRR: 53 dB
** VoutMax: 4.25 V
** VoutMin: 0.420001 V
** VcmMax: 4.24001 V
** VcmMin: 1.84001 V


** Expected Currents: 
** NormalTransistorNmos: 1.15471e+07 muA
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -1.4574e+08 muA
** DiodeTransistorPmos: -2.06641e+08 muA
** DiodeTransistorPmos: -2.06641e+08 muA
** NormalTransistorNmos: 4.13282e+08 muA
** NormalTransistorNmos: 4.13281e+08 muA
** NormalTransistorNmos: 2.06642e+08 muA
** NormalTransistorNmos: 2.06642e+08 muA
** NormalTransistorNmos: 1.92347e+08 muA
** NormalTransistorNmos: 1.92346e+08 muA
** NormalTransistorPmos: -1.92346e+08 muA
** NormalTransistorPmos: -1.92345e+08 muA
** NormalTransistorNmos: 1.92347e+08 muA
** NormalTransistorNmos: 1.92346e+08 muA
** NormalTransistorPmos: -1.92346e+08 muA
** NormalTransistorPmos: -1.92345e+08 muA
** DiodeTransistorNmos: 1.45741e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.15479e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 0.618001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.822001  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.646001  V
** out: 2.5  V
** outFirstStage: 3.83601  V
** outVoltageBiasXXpXX0: 3.76001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.213001  V
** sourceTransconductance: 1.48001  V
** innerStageBias: 0.241001  V
** innerTransconductance: 4.40001  V
** inner: 0.241001  V
** inner: 4.40001  V


.END