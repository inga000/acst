.suckt  two_stage_single_output_op_amp_140_4 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias2 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mMainBias3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad6 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
mSimpleFirstStageLoad11 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1Transconductor15 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias17 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mSecondStage1StageBias18 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos
mMainBias19 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias20 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias21 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mMainBias22 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_140_4

