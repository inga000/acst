.suckt  symmetrical_op_amp1 ibias in1 in2 out sourceNmos sourcePmos
m1 outFirstStage outFirstStage sourceNmos sourceNmos nmos
m2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m3 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m4 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m5 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c1 out sourceNmos 
m6 out outFirstStage sourceNmos sourceNmos nmos
m7 out innerComplementarySecondStage sourcePmos sourcePmos pmos
m8 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos
m9 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m10 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp1

