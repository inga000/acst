** Name: one_stage_single_output_op_amp102

.MACRO one_stage_single_output_op_amp102 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=32e-6
mMainBias2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mMainBias3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=25e-6
mTelescopicFirstStageStageBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=342e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=7e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=32e-6
mTelescopicFirstStageLoad7 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=16e-6
mMainBias8 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=27e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=52e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=104e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=104e-6
mMainBias12 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=25e-6
mMainBias13 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=12e-6
mTelescopicFirstStageLoad14 out outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=52e-6
mTelescopicFirstStageStageBias15 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=342e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp102

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 0.820001 mW
** Area: 3882 (mu_m)^2
** Transit frequency: 2.57601 MHz
** Transit frequency with error factor: 2.57637 MHz
** Slew rate: 6.94852 V/mu_s
** Phase margin: 86.5167°
** CMRR: 135 dB
** VoutMax: 3.07001 V
** VoutMin: 0.900001 V
** VcmMax: 3 V
** VcmMin: 0.830001 V


** Expected Currents: 
** NormalTransistorNmos: 2.60871e+07 muA
** NormalTransistorPmos: -4.87799e+06 muA
** NormalTransistorPmos: -5.65089e+07 muA
** NormalTransistorPmos: -5.65099e+07 muA
** NormalTransistorNmos: 5.65081e+07 muA
** NormalTransistorNmos: 5.65091e+07 muA
** DiodeTransistorNmos: 5.65081e+07 muA
** NormalTransistorPmos: -1.39104e+08 muA
** DiodeTransistorPmos: -1.39103e+08 muA
** NormalTransistorPmos: -5.65089e+07 muA
** NormalTransistorPmos: -5.65089e+07 muA
** DiodeTransistorNmos: 4.87701e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -2.60879e+07 muA


** Expected Voltages: 
** ibias: 3.35001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.590001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.17601  V
** outVoltageBiasXXpXX2: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.41101  V
** innerSourceLoad2: 0.693001  V
** out1: 1.30201  V
** sourceGCC1: 2.99401  V
** sourceGCC2: 2.99401  V
** inner: 4.17201  V


.END