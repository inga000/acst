** Name: one_stage_single_output_op_amp80

.MACRO one_stage_single_output_op_amp80 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=5e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=27e-6
m3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=24e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m6 out outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=352e-6
m7 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=144e-6
m8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=144e-6
m9 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=6e-6 W=352e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=32e-6
m11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=32e-6
m12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=27e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
m14 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=244e-6
m15 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
m16 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
m17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=244e-6
m18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=203e-6
m19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=203e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp80

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 2.41701 mW
** Area: 6077 (mu_m)^2
** Transit frequency: 6.81501 MHz
** Transit frequency with error factor: 6.81493 MHz
** Slew rate: 6.81439 V/mu_s
** Phase margin: 87.6626°
** CMRR: 147 dB
** VoutMax: 4.02001 V
** VoutMin: 0.320001 V
** VcmMax: 5.17001 V
** VcmMin: 1.81001 V


** Expected Currents: 
** NormalTransistorPmos: -2.53459e+07 muA
** NormalTransistorPmos: -2.63599e+07 muA
** NormalTransistorPmos: -1.3721e+08 muA
** NormalTransistorPmos: -2.05814e+08 muA
** NormalTransistorPmos: -1.37212e+08 muA
** NormalTransistorPmos: -2.05816e+08 muA
** NormalTransistorNmos: 1.37211e+08 muA
** NormalTransistorNmos: 1.37212e+08 muA
** NormalTransistorNmos: 1.37213e+08 muA
** NormalTransistorNmos: 1.37212e+08 muA
** NormalTransistorNmos: 1.3721e+08 muA
** DiodeTransistorNmos: 1.37209e+08 muA
** NormalTransistorNmos: 6.86051e+07 muA
** NormalTransistorNmos: 6.86051e+07 muA
** DiodeTransistorNmos: 2.53451e+07 muA
** NormalTransistorNmos: 2.53441e+07 muA
** DiodeTransistorNmos: 2.63591e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.48201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outInputVoltageBiasXXnXX1: 1.65601  V
** outSourceVoltageBiasXXnXX1: 0.828001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.921001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.349001  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.22301  V
** sourceGCC2: 4.22301  V
** sourceTransconductance: 1.93601  V
** inner: 0.826001  V


.END