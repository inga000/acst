** Name: two_stage_single_output_op_amp_75_3

.MACRO two_stage_single_output_op_amp_75_3 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=80e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=27e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=34e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=15e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=74e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=80e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=48e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=48e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=355e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=505e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=267e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=390e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=243e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=243e-6
mSecondStage1StageBias16 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=433e-6
mMainBias17 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=153e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=80e-6
mSecondStage1StageBias19 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=407e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=390e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.90001e-12
.EOM two_stage_single_output_op_amp_75_3

** Expected Performance Values: 
** Gain: 133 dB
** Power consumption: 5.94001 mW
** Area: 7511 (mu_m)^2
** Transit frequency: 8.32301 MHz
** Transit frequency with error factor: 8.32304 MHz
** Slew rate: 15.6238 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 3.95001 V
** VoutMin: 0.170001 V
** VcmMax: 5.17001 V
** VcmMin: 1.55001 V


** Expected Currents: 
** NormalTransistorPmos: -1.55122e+08 muA
** NormalTransistorPmos: -8.10789e+07 muA
** NormalTransistorPmos: -1.58392e+08 muA
** NormalTransistorPmos: -2.46371e+08 muA
** NormalTransistorPmos: -1.58392e+08 muA
** NormalTransistorPmos: -2.46371e+08 muA
** DiodeTransistorNmos: 1.58393e+08 muA
** NormalTransistorNmos: 1.58393e+08 muA
** NormalTransistorNmos: 1.58393e+08 muA
** NormalTransistorNmos: 1.75956e+08 muA
** NormalTransistorNmos: 1.75955e+08 muA
** NormalTransistorNmos: 8.79781e+07 muA
** NormalTransistorNmos: 8.79781e+07 muA
** NormalTransistorNmos: 4.3901e+08 muA
** NormalTransistorPmos: -4.39009e+08 muA
** NormalTransistorPmos: -4.39008e+08 muA
** DiodeTransistorNmos: 1.55123e+08 muA
** DiodeTransistorNmos: 8.10781e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.44101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.925001  V
** inputVoltageBiasXXnXX2: 0.572001  V
** out: 2.5  V
** outFirstStage: 0.580001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.367001  V
** innerTransistorStack2Load2: 0.353001  V
** out1: 0.558001  V
** sourceGCC1: 4.15501  V
** sourceGCC2: 4.15501  V
** sourceTransconductance: 1.67701  V
** innerStageBias: 4.25  V


.END