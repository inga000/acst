.suckt  complementary_op_amp34 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m3 FirstStageYinnerOutputLoadNmos outInputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m4 FirstStageYinnerTransistorStack1LoadPmos outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m5 out outInputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m6 FirstStageYinnerTransistorStack2LoadPmos outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m7 FirstStageYinnerOutputLoadNmos FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m8 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack2LoadNmos sourceNmos sourceNmos nmos
m9 out FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m10 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos sourceNmos sourceNmos nmos
m11 FirstStageYsourceTransconductanceNmos ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m12 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m13 FirstStageYsourceTransconductancePmos outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m14 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m15 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m16 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m17 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m18 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c1 out sourceNmos 
m19 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m20 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m21 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m23 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m24 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end complementary_op_amp34

