.suckt  symmetrical_op_amp98 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage ibias sourcePmos sourcePmos pmos
m2 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m3 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos
m4 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m5 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m6 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m7 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c1 out sourceNmos 
m9 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m10 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m11 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos
m12 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m13 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
m14 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m15 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m17 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos
m18 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp98

