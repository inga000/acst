** Name: one_stage_single_output_op_amp120

.MACRO one_stage_single_output_op_amp120 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=10e-6
mTelescopicFirstStageStageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=85e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=22e-6
mTelescopicFirstStageLoad4 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mTelescopicFirstStageLoad5 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=58e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mTelescopicFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=65e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=65e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=65e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias11 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mTelescopicFirstStageLoad12 out outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=65e-6
mTelescopicFirstStageStageBias13 sourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=85e-6
mTelescopicFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mTelescopicFirstStageLoad15 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=58e-6
mMainBias16 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=25e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp120

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 0.501001 mW
** Area: 2034 (mu_m)^2
** Transit frequency: 2.62201 MHz
** Transit frequency with error factor: 2.62213 MHz
** Slew rate: 4.16108 V/mu_s
** Phase margin: 85.9437°
** CMRR: 152 dB
** VoutMax: 4.06001 V
** VoutMin: 1.01001 V
** VcmMax: 3.75 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 6.89701e+06 muA
** NormalTransistorPmos: -3.38599e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** DiodeTransistorPmos: -2.47619e+07 muA
** DiodeTransistorPmos: -2.47629e+07 muA
** NormalTransistorPmos: -2.47619e+07 muA
** NormalTransistorPmos: -2.47629e+07 muA
** NormalTransistorNmos: 8.33821e+07 muA
** DiodeTransistorNmos: 8.33831e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 3.38591e+07 muA
** DiodeTransistorPmos: -6.89799e+06 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.04501  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.20901  V
** innerTransistorStack2Load2: 4.20801  V
** out1: 3.49001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.556001  V


.END