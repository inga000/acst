** Name: two_stage_single_output_op_amp_106_1

.MACRO two_stage_single_output_op_amp_106_1 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=21e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=378e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=18e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=5e-6
mTelescopicFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=234e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=45e-6
mTelescopicFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=273e-6
mTelescopicFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=21e-6
mMainBias11 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
mMainBias12 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=362e-6
mTelescopicFirstStageLoad13 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=34e-6
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=112e-6
mTelescopicFirstStageTransconductor15 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=7e-6 W=112e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=5e-6
mMainBias17 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=129e-6
mSecondStage1StageBias18 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=528e-6
mTelescopicFirstStageLoad19 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=34e-6
mTelescopicFirstStageStageBias20 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=234e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_106_1

** Expected Performance Values: 
** Gain: 141 dB
** Power consumption: 2.40501 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 3.76901 MHz
** Transit frequency with error factor: 3.76881 MHz
** Slew rate: 12.0622 V/mu_s
** Phase margin: 61.8795°
** CMRR: 139 dB
** VoutMax: 4.69001 V
** VoutMin: 0.300001 V
** VcmMax: 3.18001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorNmos: 1.90501e+06 muA
** NormalTransistorNmos: 6.96431e+07 muA
** NormalTransistorPmos: -7.19959e+07 muA
** NormalTransistorPmos: -1.00009e+07 muA
** NormalTransistorPmos: -1.00009e+07 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** NormalTransistorNmos: 1.00001e+07 muA
** NormalTransistorNmos: 1.00001e+07 muA
** NormalTransistorPmos: -8.96489e+07 muA
** DiodeTransistorPmos: -8.96499e+07 muA
** NormalTransistorPmos: -1.00019e+07 muA
** NormalTransistorPmos: -1.00019e+07 muA
** NormalTransistorNmos: 2.97471e+08 muA
** NormalTransistorPmos: -2.9747e+08 muA
** DiodeTransistorNmos: 7.19951e+07 muA
** DiodeTransistorPmos: -1.90599e+06 muA
** NormalTransistorPmos: -1.90699e+06 muA
** DiodeTransistorPmos: -6.96439e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outInputVoltageBiasXXpXX1: 3.36401  V
** outSourceVoltageBiasXXpXX1: 4.18201  V
** outVoltageBiasXXpXX2: 2.27201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.25101  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 3.01801  V
** sourceGCC2: 3.01701  V
** inner: 4.18001  V


.END