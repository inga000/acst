** Name: two_stage_single_output_op_amp_25_3

.MACRO two_stage_single_output_op_amp_25_3 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=52e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=52e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=52e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=241e-6
mSimpleFirstStageLoad7 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=52e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=370e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=36e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=443e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=370e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9e-12
.EOM two_stage_single_output_op_amp_25_3

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 3.41101 mW
** Area: 10070 (mu_m)^2
** Transit frequency: 5.44501 MHz
** Transit frequency with error factor: 5.43973 MHz
** Slew rate: 7.24563 V/mu_s
** Phase margin: 60.1606°
** CMRR: 102 dB
** negPSRR: 97 dB
** posPSRR: 101 dB
** VoutMax: 3.93001 V
** VoutMin: 0.380001 V
** VcmMax: 3.11001 V
** VcmMin: 0.630001 V


** Expected Currents: 
** DiodeTransistorNmos: 3.29511e+07 muA
** NormalTransistorNmos: 3.29501e+07 muA
** NormalTransistorNmos: 3.29511e+07 muA
** DiodeTransistorNmos: 3.29501e+07 muA
** NormalTransistorPmos: -6.59029e+07 muA
** NormalTransistorPmos: -6.59019e+07 muA
** NormalTransistorPmos: -3.29519e+07 muA
** NormalTransistorPmos: -3.29519e+07 muA
** NormalTransistorNmos: 5.96281e+08 muA
** NormalTransistorPmos: -5.9628e+08 muA
** NormalTransistorPmos: -5.96281e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.789001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.616001  V
** innerStageBias: 4.29201  V
** innerTransistorStack1Load1: 0.616001  V
** out1: 1.19401  V
** sourceTransconductance: 3.27501  V
** innerStageBias: 4.24701  V


.END