** Name: symmetrical_op_amp28

.MACRO symmetrical_op_amp28 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mSecondStage1StageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=24e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=6e-6 W=24e-6
mSecondStage1StageBias4 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSymmetricalFirstStageLoad5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=127e-6
mSymmetricalFirstStageLoad6 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=127e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=166e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias8 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=24e-6
mMainBias9 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos4 L=3e-6 W=68e-6
mSymmetricalFirstStageTransconductor10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=35e-6
mSecondStage1StageBias11 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=6e-6 W=24e-6
mSymmetricalFirstStageTransconductor12 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=35e-6
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=154e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor14 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=154e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=412e-6
mSecondStage1Transconductor16 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=412e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp28

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 3.65201 mW
** Area: 5923 (mu_m)^2
** Transit frequency: 5.00601 MHz
** Transit frequency with error factor: 5.00601 MHz
** Slew rate: 16.6006 V/mu_s
** Phase margin: 62.4525°
** CMRR: 126 dB
** negPSRR: 46 dB
** posPSRR: 54 dB
** VoutMax: 4.25 V
** VoutMin: 1.80001 V
** VcmMax: 4.24001 V
** VcmMin: 1.18001 V


** Expected Currents: 
** NormalTransistorNmos: 1.11687e+08 muA
** DiodeTransistorPmos: -1.37543e+08 muA
** DiodeTransistorPmos: -1.37543e+08 muA
** NormalTransistorNmos: 2.75086e+08 muA
** NormalTransistorNmos: 1.37544e+08 muA
** NormalTransistorNmos: 1.37544e+08 muA
** NormalTransistorNmos: 1.66787e+08 muA
** DiodeTransistorNmos: 1.66786e+08 muA
** NormalTransistorPmos: -1.66786e+08 muA
** NormalTransistorPmos: -1.66785e+08 muA
** DiodeTransistorNmos: 1.66787e+08 muA
** NormalTransistorNmos: 1.66786e+08 muA
** NormalTransistorPmos: -1.66786e+08 muA
** NormalTransistorPmos: -1.66785e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.11686e+08 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceStageBiasComplementarySecondStage: 1.10401  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 2.20801  V
** out: 2.5  V
** outFirstStage: 3.83601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.56501  V
** innerTransconductance: 4.40001  V
** inner: 1.09801  V
** inner: 4.40001  V


.END