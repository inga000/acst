** Name: two_stage_single_output_op_amp_78_7

.MACRO two_stage_single_output_op_amp_78_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=10e-6 W=49e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=10e-6 W=53e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=16e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=43e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=36e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=24e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=10e-6 W=49e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=23e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=23e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=43e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=16e-6
mSecondStage1StageBias13 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=467e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=53e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=182e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=83e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=83e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=348e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=182e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=24e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=283e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5e-12
.EOM two_stage_single_output_op_amp_78_7

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 10.0811 mW
** Area: 6659 (mu_m)^2
** Transit frequency: 5.48101 MHz
** Transit frequency with error factor: 5.48066 MHz
** Slew rate: 4.86211 V/mu_s
** Phase margin: 60.1606°
** CMRR: 142 dB
** VoutMax: 4.25 V
** VoutMin: 0.210001 V
** VcmMax: 5.12001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorPmos: -1.16469e+07 muA
** NormalTransistorPmos: -1.37337e+08 muA
** NormalTransistorPmos: -2.46379e+07 muA
** NormalTransistorPmos: -4.02789e+07 muA
** NormalTransistorPmos: -2.46379e+07 muA
** NormalTransistorPmos: -4.02789e+07 muA
** DiodeTransistorNmos: 2.46371e+07 muA
** DiodeTransistorNmos: 2.46361e+07 muA
** NormalTransistorNmos: 2.46371e+07 muA
** NormalTransistorNmos: 2.46361e+07 muA
** NormalTransistorNmos: 3.12791e+07 muA
** DiodeTransistorNmos: 3.12781e+07 muA
** NormalTransistorNmos: 1.56401e+07 muA
** NormalTransistorNmos: 1.56401e+07 muA
** NormalTransistorNmos: 1.7667e+09 muA
** NormalTransistorPmos: -1.76669e+09 muA
** DiodeTransistorNmos: 1.16461e+07 muA
** NormalTransistorNmos: 1.16451e+07 muA
** DiodeTransistorNmos: 1.37338e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.22401  V
** outSourceVoltageBiasXXnXX1: 0.612001  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** outVoltageBiasXXnXX2: 0.617001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.648001  V
** innerTransistorStack2Load2: 0.647001  V
** out1: 1.28701  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.91501  V
** inner: 0.611001  V


.END