.suckt  two_stage_single_output_op_amp_91_4 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m4 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m5 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m6 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m7 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m8 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos
m9 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m10 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos
m11 sourceTransconductance ibias sourcePmos sourcePmos pmos
m12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c2 out sourceNmos 
m14 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m15 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m16 out outVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m17 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos
m18 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m19 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m20 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
m21 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m22 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_91_4

