.suckt  two_stage_single_output_op_amp_185_3 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_2 FirstStageYinnerLoad1 FirstStageYinnerLoad1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_3 outFirstStage FirstStageYinnerLoad1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_4 FirstStageYinnerLoad1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_6 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m_SingleOutput_FirstStage_Load_7 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_StageBias_8 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_SingleOutput_FirstStage_StageBias_9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Transconductor_10 FirstStageYinnerLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_SingleOutput_FirstStage_Transconductor_11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_Transconductor_12 out outFirstStage sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_13 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m_SingleOutput_SecondStage1_StageBias_14 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_15 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_SingleOutput_MainBias_16 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_17 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_SingleOutput_MainBias_18 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_185_3

