.suckt  two_stage_single_output_op_amp_86_10 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXpXX3 ibias sourceNmos sourceNmos nmos
m4 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m5 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m6 FirstStageYout1 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos
m7 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m8 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos
m9 sourceTransconductance inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c2 out sourceNmos 
m12 out ibias sourceNmos sourceNmos nmos
m13 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m14 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
m15 ibias ibias sourceNmos sourceNmos nmos
m16 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
m17 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m18 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_86_10

