** Name: two_stage_single_output_op_amp_44_5

.MACRO two_stage_single_output_op_amp_44_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=17e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=120e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=11e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=376e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=21e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=88e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=88e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=58e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=21e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=104e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=7e-6 W=120e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=107e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=107e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=11e-6
mSecondStage1StageBias19 out inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=376e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=9e-6 W=239e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_44_5

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 3.24501 mW
** Area: 9788 (mu_m)^2
** Transit frequency: 3.54501 MHz
** Transit frequency with error factor: 3.54479 MHz
** Slew rate: 3.50938 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 3.63001 V
** VoutMin: 0.570001 V
** VcmMax: 4.09001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.59601e+07 muA
** NormalTransistorNmos: 2.84101e+07 muA
** NormalTransistorNmos: 1.59681e+07 muA
** NormalTransistorNmos: 2.40241e+07 muA
** NormalTransistorNmos: 1.59681e+07 muA
** NormalTransistorNmos: 2.40241e+07 muA
** NormalTransistorPmos: -1.59689e+07 muA
** NormalTransistorPmos: -1.59689e+07 muA
** DiodeTransistorPmos: -1.59689e+07 muA
** NormalTransistorPmos: -1.61149e+07 muA
** NormalTransistorPmos: -8.05699e+06 muA
** NormalTransistorPmos: -8.05699e+06 muA
** NormalTransistorNmos: 5.46524e+08 muA
** NormalTransistorPmos: -5.46523e+08 muA
** DiodeTransistorPmos: -5.46524e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.59609e+07 muA
** NormalTransistorPmos: -1.59619e+07 muA
** DiodeTransistorPmos: -2.84109e+07 muA


** Expected Voltages: 
** ibias: 1.18101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.06201  V
** out: 2.5  V
** outFirstStage: 0.976001  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outSourceVoltageBiasXXpXX1: 4.03101  V
** outVoltageBiasXXpXX2: 4.25301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.20701  V
** out1: 3.45901  V
** sourceGCC1: 0.524001  V
** sourceGCC2: 0.524001  V
** sourceTransconductance: 3.22301  V
** inner: 4.02701  V


.END