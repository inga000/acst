** Name: two_stage_single_output_op_amp_5_1

.MACRO two_stage_single_output_op_amp_5_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
mMainBias2 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mSimpleFirstStageLoad3 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=117e-6
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=167e-6
mSimpleFirstStageLoad7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=117e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=10e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=145e-6
mMainBias10 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mSecondStage1StageBias11 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=365e-6
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_5_1

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 1.25801 mW
** Area: 3471 (mu_m)^2
** Transit frequency: 3.04801 MHz
** Transit frequency with error factor: 3.04108 MHz
** Slew rate: 6.46538 V/mu_s
** Phase margin: 71.6198°
** CMRR: 93 dB
** negPSRR: 94 dB
** posPSRR: 223 dB
** VoutMax: 4.84001 V
** VoutMin: 0.150001 V
** VcmMax: 3.55001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -8.78499e+06 muA
** NormalTransistorNmos: 3.18491e+07 muA
** NormalTransistorNmos: 3.18481e+07 muA
** NormalTransistorNmos: 3.18471e+07 muA
** NormalTransistorNmos: 3.18481e+07 muA
** NormalTransistorPmos: -6.36949e+07 muA
** NormalTransistorPmos: -3.18479e+07 muA
** NormalTransistorPmos: -3.18479e+07 muA
** NormalTransistorNmos: 1.59093e+08 muA
** NormalTransistorPmos: -1.59092e+08 muA
** DiodeTransistorNmos: 8.78401e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.79201  V


.END