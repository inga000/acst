** Name: two_stage_single_output_op_amp_30_9

.MACRO two_stage_single_output_op_amp_30_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=377e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=76e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=271e-6
mSimpleFirstStageLoad5 FirstStageYinnerLoad1 FirstStageYinnerLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=71e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=105e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=53e-6
mSimpleFirstStageStageBias8 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=76e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=377e-6
mMainBias10 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias11 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=153e-6
mSecondStage1StageBias12 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=271e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=53e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=483e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYinnerLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=71e-6
mMainBias16 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=37e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_30_9

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 4.92701 mW
** Area: 11515 (mu_m)^2
** Transit frequency: 5.25301 MHz
** Transit frequency with error factor: 5.24906 MHz
** Slew rate: 4.95082 V/mu_s
** Phase margin: 74.4846°
** CMRR: 99 dB
** negPSRR: 162 dB
** posPSRR: 97 dB
** VoutMax: 4.75 V
** VoutMin: 0.840001 V
** VcmMax: 4.59001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 3.08016e+08 muA
** NormalTransistorPmos: -1.10152e+08 muA
** DiodeTransistorPmos: -1.12179e+07 muA
** NormalTransistorPmos: -1.12179e+07 muA
** NormalTransistorNmos: 2.24331e+07 muA
** DiodeTransistorNmos: 2.24321e+07 muA
** NormalTransistorNmos: 1.12171e+07 muA
** NormalTransistorNmos: 1.12171e+07 muA
** NormalTransistorNmos: 5.34767e+08 muA
** DiodeTransistorNmos: 5.34768e+08 muA
** NormalTransistorPmos: -5.34766e+08 muA
** DiodeTransistorNmos: 1.10153e+08 muA
** NormalTransistorNmos: 1.10153e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.08015e+08 muA


** Expected Voltages: 
** ibias: 1.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.73101  V
** out: 2.5  V
** outFirstStage: 4.18601  V
** outInputVoltageBiasXXnXX1: 1.14401  V
** outSourceVoltageBiasXXnXX1: 0.572001  V
** outSourceVoltageBiasXXnXX2: 0.622001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad1: 4.18601  V
** sourceTransconductance: 1.94501  V
** inner: 0.572001  V
** inner: 0.619001  V


.END