** Name: one_stage_single_output_op_amp53

.MACRO one_stage_single_output_op_amp53 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=129e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=12e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=47e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=434e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=434e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=453e-6
mMainBias10 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=82e-6
mFoldedCascodeFirstStageLoad11 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=129e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=599e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=409e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=409e-6
mFoldedCascodeFirstStageLoad15 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=599e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp53

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 4.83901 mW
** Area: 8774 (mu_m)^2
** Transit frequency: 18.3951 MHz
** Transit frequency with error factor: 18.3947 MHz
** Slew rate: 12.8744 V/mu_s
** Phase margin: 83.6519°
** CMRR: 143 dB
** VoutMax: 4.03001 V
** VoutMin: 0.980001 V
** VcmMax: 5.16001 V
** VcmMin: 0.730001 V


** Expected Currents: 
** NormalTransistorNmos: 6.82771e+07 muA
** NormalTransistorPmos: -2.59763e+08 muA
** NormalTransistorPmos: -4.44795e+08 muA
** NormalTransistorPmos: -2.59763e+08 muA
** NormalTransistorPmos: -4.44795e+08 muA
** DiodeTransistorNmos: 2.59764e+08 muA
** DiodeTransistorNmos: 2.59763e+08 muA
** NormalTransistorNmos: 2.59764e+08 muA
** NormalTransistorNmos: 2.59763e+08 muA
** NormalTransistorNmos: 3.70064e+08 muA
** NormalTransistorNmos: 1.85032e+08 muA
** NormalTransistorNmos: 1.85032e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.82779e+07 muA
** DiodeTransistorPmos: -6.82769e+07 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.18901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.765001  V
** innerTransistorStack2Load2: 0.764001  V
** out1: 1.38801  V
** sourceGCC1: 3.75501  V
** sourceGCC2: 3.75501  V
** sourceTransconductance: 1.93601  V


.END