** Name: two_stage_single_output_op_amp_114_9

.MACRO two_stage_single_output_op_amp_114_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=4e-6 W=16e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=107e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=203e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=521e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=22e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=20e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=35e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=20e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=20e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=20e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=107e-6
mMainBias12 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=16e-6
mMainBias13 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=18e-6
mSecondStage1StageBias14 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=521e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=20e-6
mTelescopicFirstStageStageBias16 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=203e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=378e-6
mTelescopicFirstStageLoad18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=20e-6
mMainBias19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=79e-6
mMainBias20 outVoltageBiasXXnXX3 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=104e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_114_9

** Expected Performance Values: 
** Gain: 103 dB
** Power consumption: 2.07201 mW
** Area: 11386 (mu_m)^2
** Transit frequency: 3.58501 MHz
** Transit frequency with error factor: 3.58327 MHz
** Slew rate: 10.7375 V/mu_s
** Phase margin: 68.755°
** CMRR: 95 dB
** VoutMax: 4.78001 V
** VoutMin: 0.75 V
** VcmMax: 4.48001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 1.12511e+07 muA
** NormalTransistorPmos: -2.54759e+07 muA
** NormalTransistorPmos: -3.31909e+07 muA
** NormalTransistorNmos: 7.61901e+06 muA
** NormalTransistorNmos: 7.61901e+06 muA
** DiodeTransistorPmos: -7.61999e+06 muA
** NormalTransistorPmos: -7.61999e+06 muA
** NormalTransistorNmos: 4.84271e+07 muA
** DiodeTransistorNmos: 4.84261e+07 muA
** NormalTransistorNmos: 7.61901e+06 muA
** NormalTransistorNmos: 7.61901e+06 muA
** NormalTransistorNmos: 3.1921e+08 muA
** DiodeTransistorNmos: 3.19211e+08 muA
** NormalTransistorPmos: -3.19209e+08 muA
** DiodeTransistorNmos: 2.54751e+07 muA
** NormalTransistorNmos: 2.54751e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 3.31901e+07 muA
** DiodeTransistorPmos: -1.12519e+07 muA


** Expected Voltages: 
** ibias: 1.15101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.13601  V
** out: 2.5  V
** outFirstStage: 4.21801  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.576001  V
** outVoltageBiasXXnXX3: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.22901  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.555001  V
** inner: 0.574001  V


.END