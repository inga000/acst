** Name: one_stage_single_output_op_amp109

.MACRO one_stage_single_output_op_amp109 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
m2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=37e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=37e-6
m4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=17e-6
m5 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
m6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=4e-6
m7 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=37e-6
m8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
m9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=37e-6
m10 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=35e-6
m11 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
m12 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=580e-6
m13 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=58e-6
m14 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=35e-6
m15 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=278e-6
m16 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=278e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp109

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 0.791001 mW
** Area: 5448 (mu_m)^2
** Transit frequency: 3.26801 MHz
** Transit frequency with error factor: 3.26808 MHz
** Slew rate: 5.8832 V/mu_s
** Phase margin: 87.0896°
** CMRR: 140 dB
** VoutMax: 3.07001 V
** VoutMin: 0.870001 V
** VcmMax: 3 V
** VcmMin: 1.21001 V


** Expected Currents: 
** NormalTransistorNmos: 1.57311e+07 muA
** NormalTransistorPmos: -2.03629e+07 muA
** NormalTransistorPmos: -5.10249e+07 muA
** NormalTransistorPmos: -5.10249e+07 muA
** DiodeTransistorNmos: 5.10241e+07 muA
** NormalTransistorNmos: 5.10231e+07 muA
** NormalTransistorNmos: 5.10241e+07 muA
** DiodeTransistorNmos: 5.10231e+07 muA
** NormalTransistorPmos: -1.17778e+08 muA
** NormalTransistorPmos: -1.17779e+08 muA
** NormalTransistorPmos: -5.10239e+07 muA
** NormalTransistorPmos: -5.10239e+07 muA
** DiodeTransistorNmos: 2.03621e+07 muA
** DiodeTransistorPmos: -1.57319e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.14001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX2: 3.96101  V
** outVoltageBiasXXnXX0: 0.636001  V
** outVoltageBiasXXpXX1: 1.93801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.31101  V
** innerSourceLoad2: 0.689001  V
** innerStageBias: 3.85401  V
** innerTransistorStack1Load2: 0.688001  V
** out1: 1.27401  V
** sourceGCC1: 2.99901  V
** sourceGCC2: 2.99601  V


.END