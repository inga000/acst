.suckt  two_stage_single_output_op_amp_143_7 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad3 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad5 FirstStageYout1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad6 outFirstStage inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSimpleFirstStageTransconductor9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias10 out ibias sourceNmos sourceNmos nmos
mSecondStage1Transconductor11 out outFirstStage sourcePmos sourcePmos pmos
mMainBias12 ibias ibias sourceNmos sourceNmos nmos
mMainBias13 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_143_7

