** Name: two_stage_single_output_op_amp_122_7

.MACRO two_stage_single_output_op_amp_122_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=58e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=123e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=5e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=23e-6
mMainBias6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=67e-6
mTelescopicFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=99e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=20e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=1e-6 W=20e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=58e-6
mMainBias11 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=37e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mTelescopicFirstStageLoad13 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=99e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=93e-6
mTelescopicFirstStageStageBias15 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=123e-6
mTelescopicFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=294e-6
mTelescopicFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=6e-6 W=294e-6
mTelescopicFirstStageLoad18 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=6e-6 W=50e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=542e-6
mTelescopicFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=50e-6
mMainBias21 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=26e-6
mMainBias22 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=5e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 19.2001e-12
.EOM two_stage_single_output_op_amp_122_7

** Expected Performance Values: 
** Gain: 137 dB
** Power consumption: 4.73901 mW
** Area: 9656 (mu_m)^2
** Transit frequency: 4.20201 MHz
** Transit frequency with error factor: 4.20189 MHz
** Slew rate: 4.35232 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.74001 V
** VoutMin: 0.200001 V
** VcmMax: 5.05001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 1.03138e+08 muA
** NormalTransistorNmos: 4.13431e+07 muA
** NormalTransistorPmos: -3.97169e+07 muA
** NormalTransistorPmos: -7.54499e+06 muA
** NormalTransistorNmos: 3.80921e+07 muA
** NormalTransistorNmos: 3.80921e+07 muA
** NormalTransistorPmos: -3.80929e+07 muA
** NormalTransistorPmos: -3.80939e+07 muA
** NormalTransistorPmos: -3.80929e+07 muA
** NormalTransistorPmos: -3.80939e+07 muA
** NormalTransistorNmos: 8.37291e+07 muA
** DiodeTransistorNmos: 8.37281e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorNmos: 6.69857e+08 muA
** NormalTransistorPmos: -6.69856e+08 muA
** DiodeTransistorNmos: 3.97161e+07 muA
** NormalTransistorNmos: 3.97151e+07 muA
** DiodeTransistorNmos: 7.54401e+06 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.03137e+08 muA
** DiodeTransistorPmos: -4.13439e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.66301  V
** out: 2.5  V
** outFirstStage: 4.17201  V
** outInputVoltageBiasXXnXX1: 1.12001  V
** outSourceVoltageBiasXXnXX1: 0.560001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 3.78301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.73101  V
** innerTransistorStack2Load2: 4.73101  V
** out1: 4.22701  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.559001  V


.END