** Name: two_stage_single_output_op_amp_30_8

.MACRO two_stage_single_output_op_amp_30_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=5e-6 W=6e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=28e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=64e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=188e-6
m6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=5e-6
m7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=34e-6
m8 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=64e-6
m9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
m10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=28e-6
m11 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=31e-6
m12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=5e-6 W=92e-6
m13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=34e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=502e-6
m15 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=188e-6
m16 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=8e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_30_8

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 1.57201 mW
** Area: 6760 (mu_m)^2
** Transit frequency: 5.00101 MHz
** Transit frequency with error factor: 4.99471 MHz
** Slew rate: 4.71329 V/mu_s
** Phase margin: 60.1606°
** CMRR: 102 dB
** negPSRR: 165 dB
** posPSRR: 101 dB
** VoutMax: 4.84001 V
** VoutMin: 0.940001 V
** VcmMax: 4.68001 V
** VcmMin: 1.32001 V


** Expected Currents: 
** NormalTransistorNmos: 1.18251e+07 muA
** NormalTransistorPmos: -1.85909e+07 muA
** DiodeTransistorPmos: -2.15869e+07 muA
** NormalTransistorPmos: -2.15869e+07 muA
** NormalTransistorNmos: 4.31711e+07 muA
** DiodeTransistorNmos: 4.31701e+07 muA
** NormalTransistorNmos: 2.15861e+07 muA
** NormalTransistorNmos: 2.15861e+07 muA
** NormalTransistorNmos: 2.30865e+08 muA
** NormalTransistorNmos: 2.30864e+08 muA
** NormalTransistorPmos: -2.30864e+08 muA
** DiodeTransistorNmos: 1.85901e+07 muA
** NormalTransistorNmos: 1.85891e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.18259e+07 muA


** Expected Voltages: 
** ibias: 1.27301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.80901  V
** out: 2.5  V
** outFirstStage: 4.27501  V
** outInputVoltageBiasXXnXX1: 1.16601  V
** outSourceVoltageBiasXXnXX1: 0.583001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.27501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.482001  V
** inner: 0.583001  V


.END