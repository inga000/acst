** Name: two_stage_single_output_op_amp_3_1

.MACRO two_stage_single_output_op_amp_3_1 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=53e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=17e-6
m4 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=38e-6
m5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=53e-6
m6 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=119e-6
m7 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=38e-6
m8 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=171e-6
m9 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=40e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=40e-6
m11 out ibias sourcePmos sourcePmos pmos4 L=4e-6 W=192e-6
Capacitor1 outFirstStage out 7.10001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_3_1

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 1.29101 mW
** Area: 2848 (mu_m)^2
** Transit frequency: 3.01001 MHz
** Transit frequency with error factor: 2.99897 MHz
** Slew rate: 4.19637 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** negPSRR: 94 dB
** posPSRR: 202 dB
** VoutMax: 4.64001 V
** VoutMin: 0.150001 V
** VcmMax: 3.32001 V
** VcmMin: 0.170001 V


** Expected Currents: 
** NormalTransistorPmos: -2.27199e+07 muA
** DiodeTransistorNmos: 5.07681e+07 muA
** NormalTransistorNmos: 5.07671e+07 muA
** NormalTransistorNmos: 5.07681e+07 muA
** NormalTransistorPmos: -1.01534e+08 muA
** NormalTransistorPmos: -5.07669e+07 muA
** NormalTransistorPmos: -5.07669e+07 muA
** NormalTransistorNmos: 1.13986e+08 muA
** NormalTransistorPmos: -1.13985e+08 muA
** DiodeTransistorNmos: 2.27191e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.07201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.732001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.81401  V


.END