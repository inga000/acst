** Name: two_stage_single_output_op_amp_62_10

.MACRO two_stage_single_output_op_amp_62_10 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=9e-6
m2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=116e-6
m3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=13e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=141e-6
m6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=341e-6
m7 inputVoltageBiasXXpXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=79e-6
m8 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=581e-6
m9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=54e-6
m10 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=54e-6
m11 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=69e-6
m12 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=69e-6
m13 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=79e-6
m14 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=284e-6
m15 out inputVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=592e-6
m16 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=86e-6
m17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=341e-6
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=452e-6
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=452e-6
m20 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=141e-6
m21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=13e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 8.10001e-12
.EOM two_stage_single_output_op_amp_62_10

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 9.12601 mW
** Area: 14996 (mu_m)^2
** Transit frequency: 8.69101 MHz
** Transit frequency with error factor: 8.69133 MHz
** Slew rate: 9.46306 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 4.36001 V
** VoutMin: 0.150001 V
** VcmMax: 3.04001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.51986e+08 muA
** NormalTransistorPmos: -6.16009e+07 muA
** NormalTransistorPmos: -2.20937e+08 muA
** NormalTransistorNmos: 7.69971e+07 muA
** NormalTransistorNmos: 1.31997e+08 muA
** NormalTransistorNmos: 7.69941e+07 muA
** NormalTransistorNmos: 1.31992e+08 muA
** DiodeTransistorPmos: -7.69959e+07 muA
** NormalTransistorPmos: -7.69949e+07 muA
** NormalTransistorPmos: -7.69959e+07 muA
** NormalTransistorPmos: -1.09995e+08 muA
** DiodeTransistorPmos: -1.09994e+08 muA
** NormalTransistorPmos: -5.49979e+07 muA
** NormalTransistorPmos: -5.49979e+07 muA
** NormalTransistorNmos: 1.10659e+09 muA
** NormalTransistorPmos: -1.10658e+09 muA
** NormalTransistorPmos: -1.10658e+09 muA
** DiodeTransistorNmos: 6.16001e+07 muA
** DiodeTransistorNmos: 2.20938e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -1.51985e+08 muA


** Expected Voltages: 
** ibias: 3.28201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.04401  V
** inputVoltageBiasXXnXX2: 0.555001  V
** inputVoltageBiasXXpXX2: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.11301  V
** outSourceVoltageBiasXXpXX1: 4.14201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.47301  V
** out1: 4.21101  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.31101  V
** innerTransconductance: 4.57201  V
** inner: 4.13801  V


.END