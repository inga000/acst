** Name: two_stage_single_output_op_amp_108_2

.MACRO two_stage_single_output_op_amp_108_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=25e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=171e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=16e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=8e-6
mTelescopicFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=211e-6
mTelescopicFirstStageLoad7 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=35e-6
mTelescopicFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=78e-6
mTelescopicFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=78e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=494e-6
mMainBias11 inputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=191e-6
mSecondStage1Transconductor12 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=394e-6
mTelescopicFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=35e-6
mMainBias14 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=14e-6
mTelescopicFirstStageLoad15 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=6e-6 W=17e-6
mTelescopicFirstStageTransconductor16 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=177e-6
mTelescopicFirstStageTransconductor17 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=177e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
mMainBias19 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=109e-6
mSecondStage1StageBias20 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=438e-6
mTelescopicFirstStageLoad21 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=6e-6 W=17e-6
mMainBias22 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=75e-6
mTelescopicFirstStageStageBias23 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=211e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.30001e-12
.EOM two_stage_single_output_op_amp_108_2

** Expected Performance Values: 
** Gain: 143 dB
** Power consumption: 1.81001 mW
** Area: 14951 (mu_m)^2
** Transit frequency: 2.77901 MHz
** Transit frequency with error factor: 2.77882 MHz
** Slew rate: 6.65551 V/mu_s
** Phase margin: 60.1606°
** CMRR: 136 dB
** VoutMax: 4.84001 V
** VoutMin: 0.300001 V
** VcmMax: 3.26001 V
** VcmMin: 0.160001 V


** Expected Currents: 
** NormalTransistorNmos: 2.66701e+06 muA
** NormalTransistorNmos: 3.66831e+07 muA
** NormalTransistorPmos: -3.25709e+07 muA
** NormalTransistorPmos: -4.71459e+07 muA
** NormalTransistorPmos: -1.66669e+07 muA
** NormalTransistorPmos: -1.66669e+07 muA
** NormalTransistorNmos: 1.66661e+07 muA
** NormalTransistorNmos: 1.66651e+07 muA
** NormalTransistorNmos: 1.66661e+07 muA
** NormalTransistorNmos: 1.66651e+07 muA
** NormalTransistorPmos: -7.00209e+07 muA
** DiodeTransistorPmos: -7.00219e+07 muA
** NormalTransistorPmos: -1.66679e+07 muA
** NormalTransistorPmos: -1.66679e+07 muA
** NormalTransistorNmos: 1.89501e+08 muA
** NormalTransistorNmos: 1.895e+08 muA
** NormalTransistorPmos: -1.895e+08 muA
** DiodeTransistorNmos: 3.25701e+07 muA
** DiodeTransistorNmos: 4.71451e+07 muA
** DiodeTransistorPmos: -2.66799e+06 muA
** NormalTransistorPmos: -2.66899e+06 muA
** DiodeTransistorPmos: -3.66839e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXpXX2: 1.85601  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.48601  V
** outSourceVoltageBiasXXpXX1: 4.24301  V
** outVoltageBiasXXnXX0: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.29301  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** sourceGCC1: 2.99601  V
** sourceGCC2: 2.99101  V
** innerTransconductance: 0.150001  V
** inner: 4.24301  V


.END