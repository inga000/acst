** Name: two_stage_single_output_op_amp_104_7

.MACRO two_stage_single_output_op_amp_104_7 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=134e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=55e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=73e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=11e-6
mTelescopicFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=91e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=10e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=134e-6
mSecondStage1StageBias8 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=596e-6
mTelescopicFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=120e-6
mMainBias10 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mTelescopicFirstStageLoad11 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=71e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=56e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=56e-6
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mMainBias15 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=57e-6
mMainBias16 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=262e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=293e-6
mTelescopicFirstStageLoad18 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=71e-6
mTelescopicFirstStageStageBias19 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=91e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.1001e-12
.EOM two_stage_single_output_op_amp_104_7

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 11.7721 mW
** Area: 8116 (mu_m)^2
** Transit frequency: 3.75401 MHz
** Transit frequency with error factor: 3.75392 MHz
** Slew rate: 8.26705 V/mu_s
** Phase margin: 60.1606°
** CMRR: 148 dB
** VoutMax: 3.37001 V
** VoutMin: 0.280001 V
** VcmMax: 3.18001 V
** VcmMin: 0.290001 V


** Expected Currents: 
** NormalTransistorNmos: 2.66421e+07 muA
** NormalTransistorPmos: -5.25509e+07 muA
** NormalTransistorPmos: -2.39837e+08 muA
** NormalTransistorPmos: -2.86289e+07 muA
** NormalTransistorPmos: -2.86279e+07 muA
** DiodeTransistorNmos: 2.86281e+07 muA
** NormalTransistorNmos: 2.86271e+07 muA
** NormalTransistorNmos: 2.86281e+07 muA
** NormalTransistorPmos: -8.38979e+07 muA
** DiodeTransistorPmos: -8.38969e+07 muA
** NormalTransistorPmos: -2.86279e+07 muA
** NormalTransistorPmos: -2.86279e+07 muA
** NormalTransistorNmos: 1.95812e+09 muA
** NormalTransistorPmos: -1.95811e+09 muA
** DiodeTransistorNmos: 5.25501e+07 muA
** DiodeTransistorNmos: 2.39838e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -2.66429e+07 muA


** Expected Voltages: 
** ibias: 3.41801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** inputVoltageBiasXXnXX2: 0.685001  V
** out: 2.5  V
** outFirstStage: 2.81001  V
** outSourceVoltageBiasXXpXX1: 4.21001  V
** outVoltageBiasXXpXX2: 2.35001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.30201  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.06401  V
** sourceGCC2: 3.06401  V
** inner: 4.20701  V


.END