** Name: two_stage_single_output_op_amp_64_7

.MACRO two_stage_single_output_op_amp_64_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=32e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=56e-6
m3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=19e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=41e-6
m5 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=32e-6
m6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
m7 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=554e-6
m8 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=9e-6 W=42e-6
m9 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=9e-6 W=42e-6
m10 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=17e-6
m11 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=17e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=211e-6
m13 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=32e-6
m14 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=190e-6
m15 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=201e-6
m16 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=72e-6
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=72e-6
m19 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=41e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_64_7

** Expected Performance Values: 
** Gain: 117 dB
** Power consumption: 6.73801 mW
** Area: 4607 (mu_m)^2
** Transit frequency: 3.41501 MHz
** Transit frequency with error factor: 3.4149 MHz
** Slew rate: 4.74235 V/mu_s
** Phase margin: 64.1713°
** CMRR: 140 dB
** VoutMax: 4.25 V
** VoutMin: 0.150001 V
** VcmMax: 3.05001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.0094e+08 muA
** NormalTransistorPmos: -1.0666e+08 muA
** NormalTransistorNmos: 2.14241e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 2.14241e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** DiodeTransistorPmos: -2.14249e+07 muA
** DiodeTransistorPmos: -2.14259e+07 muA
** NormalTransistorPmos: -2.14249e+07 muA
** NormalTransistorPmos: -2.14259e+07 muA
** NormalTransistorPmos: -2.19079e+07 muA
** DiodeTransistorPmos: -2.19069e+07 muA
** NormalTransistorPmos: -1.09539e+07 muA
** NormalTransistorPmos: -1.09539e+07 muA
** NormalTransistorNmos: 1.05517e+09 muA
** NormalTransistorPmos: -1.05516e+09 muA
** DiodeTransistorNmos: 1.00941e+08 muA
** DiodeTransistorNmos: 1.06661e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.27301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.13801  V
** outVoltageBiasXXnXX1: 0.987001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 3.41901  V
** innerTransistorStack1Load2: 4.17701  V
** innerTransistorStack2Load2: 4.17601  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.28901  V
** inner: 4.13301  V


.END