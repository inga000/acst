.suckt  symmetrical_op_amp189 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_MainBias_1 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Load_2 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m_Symmetrical_FirstStage_Load_3 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_4 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_Symmetrical_FirstStage_Load_5 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_StageBias_6 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_Symmetrical_FirstStage_StageBias_7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Transconductor_8 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_Symmetrical_FirstStage_Transconductor_9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_StageBias_10 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos
m_Symmetrical_SecondStage1_StageBias_11 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_Transconductor_12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m_Symmetrical_SecondStage1_Transconductor_13 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_14 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_15 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_16 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_MainBias_18 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_Symmetrical_MainBias_19 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_20 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos
.end symmetrical_op_amp189

