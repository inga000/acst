** Name: two_stage_single_output_op_amp_47_7

.MACRO two_stage_single_output_op_amp_47_7 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=31e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=87e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
m5 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
m6 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=335e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=22e-6
m8 FirstStageYinnerSourceLoad2 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=22e-6
m9 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=130e-6
m10 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=130e-6
m11 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=475e-6
m12 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=86e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=246e-6
m14 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=349e-6
m15 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=6e-6 W=349e-6
m16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=50e-6
m17 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=50e-6
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=44e-6
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=44e-6
m20 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=298e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_47_7

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 1.39001 mW
** Area: 14982 (mu_m)^2
** Transit frequency: 2.67501 MHz
** Transit frequency with error factor: 2.67454 MHz
** Slew rate: 4.31923 V/mu_s
** Phase margin: 64.7443°
** CMRR: 137 dB
** VoutMax: 4.84001 V
** VoutMin: 0.150001 V
** VcmMax: 3.80001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.80901e+06 muA
** NormalTransistorPmos: -5.45e+07 muA
** NormalTransistorPmos: -9.84199e+06 muA
** NormalTransistorNmos: 2.40721e+07 muA
** NormalTransistorNmos: 4.12671e+07 muA
** NormalTransistorNmos: 2.40721e+07 muA
** NormalTransistorNmos: 4.12671e+07 muA
** NormalTransistorPmos: -2.40729e+07 muA
** NormalTransistorPmos: -2.40739e+07 muA
** NormalTransistorPmos: -2.40729e+07 muA
** NormalTransistorPmos: -2.40739e+07 muA
** NormalTransistorPmos: -3.43889e+07 muA
** NormalTransistorPmos: -1.71939e+07 muA
** NormalTransistorPmos: -1.71939e+07 muA
** NormalTransistorNmos: 1.06343e+08 muA
** NormalTransistorPmos: -1.06342e+08 muA
** DiodeTransistorNmos: 5.44991e+07 muA
** DiodeTransistorNmos: 9.84101e+06 muA
** DiodeTransistorPmos: -4.80999e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.23901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.915001  V
** inputVoltageBiasXXnXX2: 0.555001  V
** inputVoltageBiasXXpXX1: 3.91601  V
** out: 2.5  V
** outFirstStage: 4.28001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.27201  V
** innerTransistorStack1Load2: 4.63201  V
** innerTransistorStack2Load2: 4.63201  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.50601  V


.END