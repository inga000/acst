** Name: two_stage_single_output_op_amp_23_3

.MACRO two_stage_single_output_op_amp_23_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias2 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=19e-6
mMainBias3 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=426e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=35e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=35e-6
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=498e-6
mSimpleFirstStageLoad8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=426e-6
mSimpleFirstStageTransconductor9 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=383e-6
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=229e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=218e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=477e-6
mMainBias13 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=25e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=600e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=383e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.70001e-12
.EOM two_stage_single_output_op_amp_23_3

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 3.76201 mW
** Area: 14995 (mu_m)^2
** Transit frequency: 11.1861 MHz
** Transit frequency with error factor: 11.1664 MHz
** Slew rate: 16.4127 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** negPSRR: 100 dB
** posPSRR: 231 dB
** VoutMax: 3.99001 V
** VoutMin: 0.150001 V
** VcmMax: 3.03001 V
** VcmMin: -0.169999 V


** Expected Currents: 
** NormalTransistorPmos: -2.53049e+07 muA
** NormalTransistorNmos: 1.16092e+08 muA
** NormalTransistorNmos: 1.16091e+08 muA
** NormalTransistorNmos: 1.1609e+08 muA
** NormalTransistorNmos: 1.16091e+08 muA
** NormalTransistorPmos: -2.32178e+08 muA
** NormalTransistorPmos: -2.32177e+08 muA
** NormalTransistorPmos: -1.16089e+08 muA
** NormalTransistorPmos: -1.16089e+08 muA
** NormalTransistorNmos: 4.74979e+08 muA
** NormalTransistorPmos: -4.74978e+08 muA
** NormalTransistorPmos: -4.74979e+08 muA
** DiodeTransistorNmos: 2.53041e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.46301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.949001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.799001  V
** innerStageBias: 4.27001  V
** innerTransistorStack1Load1: 0.394001  V
** innerTransistorStack2Load1: 0.394001  V
** sourceTransconductance: 3.43101  V
** innerStageBias: 4.23701  V


.END