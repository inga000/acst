** Name: two_stage_single_output_op_amp_71_7

.MACRO two_stage_single_output_op_amp_71_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=28e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
m3 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=76e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=10e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=24e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=386e-6
m7 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=76e-6
m8 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
m9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=51e-6
m10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=51e-6
m11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=87e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=203e-6
m13 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=36e-6
m14 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=301e-6
m15 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=248e-6
m16 FirstStageYinnerLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=36e-6
m17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=165e-6
m18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=165e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 5.10001e-12
.EOM two_stage_single_output_op_amp_71_7

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 12.2701 mW
** Area: 5162 (mu_m)^2
** Transit frequency: 9.85901 MHz
** Transit frequency with error factor: 9.85 MHz
** Slew rate: 7.99026 V/mu_s
** Phase margin: 60.1606°
** CMRR: 106 dB
** VoutMax: 4.25 V
** VoutMin: 0.25 V
** VcmMax: 5.19001 V
** VcmMin: 1.52001 V


** Expected Currents: 
** NormalTransistorPmos: -1.27921e+08 muA
** NormalTransistorPmos: -1.04765e+08 muA
** NormalTransistorPmos: -4.09459e+07 muA
** NormalTransistorPmos: -7.01229e+07 muA
** NormalTransistorPmos: -4.09459e+07 muA
** NormalTransistorPmos: -7.01229e+07 muA
** DiodeTransistorNmos: 4.09451e+07 muA
** NormalTransistorNmos: 4.09451e+07 muA
** NormalTransistorNmos: 5.83511e+07 muA
** NormalTransistorNmos: 5.83501e+07 muA
** NormalTransistorNmos: 2.91761e+07 muA
** NormalTransistorNmos: 2.91761e+07 muA
** NormalTransistorNmos: 2.06115e+09 muA
** NormalTransistorPmos: -2.06114e+09 muA
** DiodeTransistorNmos: 1.27922e+08 muA
** DiodeTransistorNmos: 1.04766e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.21901  V
** outVoltageBiasXXnXX1: 1.13601  V
** outVoltageBiasXXnXX2: 0.655001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.600001  V
** innerStageBias: 0.450001  V
** sourceGCC1: 4.24101  V
** sourceGCC2: 4.24101  V
** sourceTransconductance: 1.91101  V


.END