** Name: two_stage_single_output_op_amp_59_1

.MACRO two_stage_single_output_op_amp_59_1 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=12e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=224e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=9e-6 W=15e-6
m5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=26e-6
m7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=89e-6
m8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=89e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=33e-6
m10 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=26e-6
m11 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=34e-6
m12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=37e-6
m13 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
m14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=224e-6
m15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=57e-6
m16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=57e-6
m17 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=9e-6 W=262e-6
m18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=527e-6
m19 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=32e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_59_1

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 4.79601 mW
** Area: 6470 (mu_m)^2
** Transit frequency: 6.01701 MHz
** Transit frequency with error factor: 6.0169 MHz
** Slew rate: 6.21644 V/mu_s
** Phase margin: 61.3065°
** CMRR: 141 dB
** VoutMax: 4.70001 V
** VoutMin: 0.550001 V
** VcmMax: 3.17001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.63171e+07 muA
** NormalTransistorNmos: 1.76311e+07 muA
** NormalTransistorNmos: 2.80721e+07 muA
** NormalTransistorNmos: 4.23781e+07 muA
** NormalTransistorNmos: 2.80721e+07 muA
** NormalTransistorNmos: 4.23781e+07 muA
** NormalTransistorPmos: -2.80729e+07 muA
** NormalTransistorPmos: -2.80729e+07 muA
** DiodeTransistorPmos: -2.80729e+07 muA
** NormalTransistorPmos: -2.86149e+07 muA
** NormalTransistorPmos: -2.86159e+07 muA
** NormalTransistorPmos: -1.43069e+07 muA
** NormalTransistorPmos: -1.43069e+07 muA
** NormalTransistorNmos: 8.3058e+08 muA
** NormalTransistorPmos: -8.30579e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.63179e+07 muA
** DiodeTransistorPmos: -1.76319e+07 muA


** Expected Voltages: 
** ibias: 1.15801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.953001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 3.69301  V
** outVoltageBiasXXpXX2: 4.13801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.26801  V
** innerStageBias: 4.49101  V
** out1: 3.48201  V
** sourceGCC1: 0.526001  V
** sourceGCC2: 0.526001  V
** sourceTransconductance: 3.23101  V


.END