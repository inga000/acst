** Name: two_stage_single_output_op_amp_73_10

.MACRO two_stage_single_output_op_amp_73_10 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=113e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=13e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=38e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=25e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=7e-6 W=113e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=13e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=45e-6
mSecondStage1StageBias11 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=400e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=10e-6 W=16e-6
mMainBias13 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=22e-6
mMainBias14 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=241e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=286e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=286e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mMainBias19 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=9e-6 W=213e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=582e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=241e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.9001e-12
.EOM two_stage_single_output_op_amp_73_10

** Expected Performance Values: 
** Gain: 134 dB
** Power consumption: 5.33901 mW
** Area: 14981 (mu_m)^2
** Transit frequency: 4.04801 MHz
** Transit frequency with error factor: 4.04788 MHz
** Slew rate: 3.81506 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 4.25 V
** VoutMin: 0.310001 V
** VcmMax: 5.04001 V
** VcmMin: 1.46001 V


** Expected Currents: 
** NormalTransistorNmos: 4.39971e+07 muA
** NormalTransistorNmos: 9.81001e+06 muA
** NormalTransistorPmos: -5.52289e+07 muA
** NormalTransistorPmos: -4.95229e+07 muA
** NormalTransistorPmos: -7.42829e+07 muA
** NormalTransistorPmos: -4.95259e+07 muA
** NormalTransistorPmos: -7.42879e+07 muA
** NormalTransistorNmos: 4.95241e+07 muA
** NormalTransistorNmos: 4.95251e+07 muA
** DiodeTransistorNmos: 4.95241e+07 muA
** NormalTransistorNmos: 4.95211e+07 muA
** NormalTransistorNmos: 4.95201e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 2.47611e+07 muA
** NormalTransistorNmos: 8.00104e+08 muA
** NormalTransistorPmos: -8.00103e+08 muA
** NormalTransistorPmos: -8.00104e+08 muA
** DiodeTransistorNmos: 5.52281e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -4.39979e+07 muA
** DiodeTransistorPmos: -9.81099e+06 muA


** Expected Voltages: 
** ibias: 0.711001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.10801  V
** out: 2.5  V
** outFirstStage: 4.16401  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.07401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.595001  V
** innerStageBias: 0.506001  V
** out1: 1.60201  V
** sourceGCC1: 4.43501  V
** sourceGCC2: 4.43501  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.72801  V


.END