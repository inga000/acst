** Name: two_stage_single_output_op_amp_10_8

.MACRO two_stage_single_output_op_amp_10_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=5e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=14e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=32e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=26e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=29e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=515e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=106e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=29e-6
mMainBias11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=14e-6
mMainBias14 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=98e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=265e-6
mSimpleFirstStageLoad16 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=8e-6 W=200e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_10_8

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 3.50001 mW
** Area: 5643 (mu_m)^2
** Transit frequency: 3.66001 MHz
** Transit frequency with error factor: 3.65703 MHz
** Slew rate: 4.42397 V/mu_s
** Phase margin: 65.8902°
** CMRR: 96 dB
** negPSRR: 160 dB
** posPSRR: 94 dB
** VoutMax: 4.40001 V
** VoutMin: 0.670001 V
** VcmMax: 4.09001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorNmos: 1.53971e+07 muA
** NormalTransistorNmos: 3.29971e+07 muA
** NormalTransistorPmos: -4.74079e+07 muA
** DiodeTransistorPmos: -1.00989e+07 muA
** NormalTransistorPmos: -1.00989e+07 muA
** NormalTransistorPmos: -1.00989e+07 muA
** NormalTransistorNmos: 2.01951e+07 muA
** NormalTransistorNmos: 1.00981e+07 muA
** NormalTransistorNmos: 1.00981e+07 muA
** NormalTransistorNmos: 5.74006e+08 muA
** NormalTransistorNmos: 5.74005e+08 muA
** NormalTransistorPmos: -5.74005e+08 muA
** DiodeTransistorNmos: 4.74071e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.53979e+07 muA
** DiodeTransistorPmos: -3.29979e+07 muA


** Expected Voltages: 
** ibias: 0.567001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.07101  V
** out: 2.5  V
** outFirstStage: 3.83601  V
** outVoltageBiasXXpXX0: 4.06801  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.40001  V
** out1: 3.83601  V
** sourceTransconductance: 1.90201  V
** innerStageBias: 0.162001  V


.END