.suckt  complementary_op_amp6 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 FirstStageYinnerSourceLoadPmos outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m5 FirstStageYinnerTransistorStack1LoadNmos inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m6 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m7 FirstStageYinnerTransistorStack2LoadNmos inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m8 FirstStageYinnerSourceLoadPmos outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m9 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m10 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m11 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m12 FirstStageYsourceTransconductanceNmos inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m13 FirstStageYsourceTransconductancePmos ibias sourcePmos sourcePmos pmos
m14 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m15 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m16 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m17 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c1 out sourceNmos 
m18 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m19 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m20 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m21 ibias ibias sourcePmos sourcePmos pmos
.end complementary_op_amp6

