** Name: two_stage_single_output_op_amp_33_8

.MACRO two_stage_single_output_op_amp_33_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=6e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
m4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=41e-6
m5 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m6 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=221e-6
m7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=21e-6
m8 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=21e-6
m9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=84e-6
m10 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=47e-6
m11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=346e-6
m13 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=145e-6
m14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=41e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_33_8

** Expected Performance Values: 
** Gain: 105 dB
** Power consumption: 1.74301 mW
** Area: 5354 (mu_m)^2
** Transit frequency: 4.63701 MHz
** Transit frequency with error factor: 4.63413 MHz
** Slew rate: 4.37002 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** negPSRR: 121 dB
** posPSRR: 105 dB
** VoutMax: 4.78001 V
** VoutMin: 0.800001 V
** VcmMax: 4.34001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2e+07 muA
** NormalTransistorPmos: -2e+07 muA
** NormalTransistorPmos: -2e+07 muA
** NormalTransistorNmos: 3.99971e+07 muA
** NormalTransistorNmos: 3.99981e+07 muA
** NormalTransistorNmos: 1.99991e+07 muA
** NormalTransistorNmos: 1.99991e+07 muA
** NormalTransistorNmos: 2.88581e+08 muA
** NormalTransistorNmos: 2.8858e+08 muA
** NormalTransistorPmos: -2.8858e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.00009e+07 muA


** Expected Voltages: 
** ibias: 1.24001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.21901  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.10601  V
** innerStageBias: 0.634001  V
** innerTransistorStack2Load1: 4.42501  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.586001  V


.END