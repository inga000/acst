.suckt  one_stage_fully_differential_op_amp9 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
m1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m3 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m4 outFeedback outFeedback sourceNmos sourceNmos nmos
m5 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m7 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m8 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m9 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m10 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m11 out1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m12 out2 outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m13 out1 outFeedback sourceNmos sourceNmos nmos
m14 out2 outFeedback sourceNmos sourceNmos nmos
m15 sourceTransconductance ibias sourcePmos sourcePmos pmos
m16 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m17 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c1 out1 sourceNmos 
c2 out2 sourceNmos 
m18 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m19 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
m20 ibias ibias sourcePmos sourcePmos pmos
.end one_stage_fully_differential_op_amp9

