** Name: two_stage_single_output_op_amp_134_3

.MACRO two_stage_single_output_op_amp_134_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=15e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mSimpleFirstStageLoad3 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=9e-6 W=27e-6
mSimpleFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=9e-6 W=27e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=224e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=122e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=122e-6
mSimpleFirstStageLoad9 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=62e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=520e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=294e-6
mSimpleFirstStageLoad12 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=62e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=458e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack1Load1 sourcePmos sourcePmos pmos4 L=9e-6 W=27e-6
mSimpleFirstStageTransconductor15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=10e-6
mSimpleFirstStageStageBias16 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=76e-6
mSecondStage1StageBias17 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSecondStage1StageBias18 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=197e-6
mSimpleFirstStageLoad19 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=9e-6 W=27e-6
mSimpleFirstStageTransconductor20 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.5e-12
.EOM two_stage_single_output_op_amp_134_3

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 8.12701 mW
** Area: 7153 (mu_m)^2
** Transit frequency: 2.51201 MHz
** Transit frequency with error factor: 2.50961 MHz
** Slew rate: 11.8974 V/mu_s
** Phase margin: 60.1606°
** CMRR: 74 dB
** VoutMax: 4.25 V
** VoutMin: 0.310001 V
** VcmMax: 3.41001 V
** VcmMin: -0.189999 V


** Expected Currents: 
** NormalTransistorNmos: 3.45215e+08 muA
** NormalTransistorNmos: 3.01344e+08 muA
** DiodeTransistorPmos: -3.04599e+07 muA
** DiodeTransistorPmos: -3.04599e+07 muA
** NormalTransistorPmos: -3.04599e+07 muA
** NormalTransistorPmos: -3.04599e+07 muA
** NormalTransistorNmos: 8.12261e+07 muA
** NormalTransistorNmos: 8.12251e+07 muA
** NormalTransistorNmos: 8.12261e+07 muA
** NormalTransistorNmos: 8.12251e+07 muA
** NormalTransistorPmos: -1.01534e+08 muA
** NormalTransistorPmos: -5.07669e+07 muA
** NormalTransistorPmos: -5.07669e+07 muA
** NormalTransistorNmos: 8.06434e+08 muA
** NormalTransistorPmos: -8.06433e+08 muA
** NormalTransistorPmos: -8.06434e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.45214e+08 muA
** DiodeTransistorPmos: -3.01343e+08 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.717001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX2: 4.16301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.495001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.495001  V
** out1: 2.37201  V
** sourceTransconductance: 3.81401  V
** innerStageBias: 4.72701  V


.END