** Name: two_stage_single_output_op_amp_30_7

.MACRO two_stage_single_output_op_amp_30_7 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=36e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=37e-6
m4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=50e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=20e-6
m6 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=18e-6
m7 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=588e-6
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=59e-6
m9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=59e-6
m10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=37e-6
m11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=36e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=97e-6
m13 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=20e-6
m14 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=74e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 8.60001e-12
.EOM two_stage_single_output_op_amp_30_7

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 5.56401 mW
** Area: 3791 (mu_m)^2
** Transit frequency: 4.68501 MHz
** Transit frequency with error factor: 4.67824 MHz
** Slew rate: 5.23496 V/mu_s
** Phase margin: 60.1606°
** CMRR: 87 dB
** negPSRR: 171 dB
** posPSRR: 86 dB
** VoutMax: 4.25 V
** VoutMin: 0.200001 V
** VcmMax: 4.09001 V
** VcmMin: 1.33001 V


** Expected Currents: 
** NormalTransistorNmos: 2.96881e+07 muA
** NormalTransistorPmos: -4.30889e+07 muA
** DiodeTransistorPmos: -2.25629e+07 muA
** NormalTransistorPmos: -2.25629e+07 muA
** NormalTransistorNmos: 4.51231e+07 muA
** DiodeTransistorNmos: 4.51221e+07 muA
** NormalTransistorNmos: 2.25621e+07 muA
** NormalTransistorNmos: 2.25621e+07 muA
** NormalTransistorNmos: 9.8488e+08 muA
** NormalTransistorPmos: -9.84879e+08 muA
** DiodeTransistorNmos: 4.30881e+07 muA
** NormalTransistorNmos: 4.30881e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.96889e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.92301  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.14801  V
** outSourceVoltageBiasXXnXX1: 0.574001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.68601  V
** sourceTransconductance: 1.91701  V
** inner: 0.574001  V


.END