.suckt  two_stage_fully_differential_op_amp_13_9 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m3 outInputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m5 outFeedback outFeedback sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m7 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m8 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m9 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m10 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m12 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m13 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m14 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m15 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m16 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m17 out1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m18 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m19 out1 out1FirstStage sourcePmos sourcePmos pmos
m20 out2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m21 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m22 out2 out2FirstStage sourcePmos sourcePmos pmos
m23 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m24 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m25 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
m26 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m27 ibias ibias sourceNmos sourceNmos nmos
m28 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_13_9

