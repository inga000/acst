.suckt  symmetrical_op_amp150 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad2 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
mSymmetricalFirstStageLoad3 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageLoad4 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
mSymmetricalFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mSymmetricalFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mSymmetricalFirstStageTransconductor8 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1Transconductor10 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mSecondStage1Transconductor11 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias12 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mSecondStage1StageBias13 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias14 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias15 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mMainBias18 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos
mMainBias19 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end symmetrical_op_amp150

