** Name: two_stage_single_output_op_amp_80_9

.MACRO two_stage_single_output_op_amp_80_9 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=13e-6
m2 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=4e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=433e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=470e-6
m5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m8 outFirstStage outVoltageBiasXXnXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=302e-6
m9 out outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=470e-6
m10 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=160e-6
m11 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=160e-6
m12 FirstStageYout1 outVoltageBiasXXnXX3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=302e-6
m13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=28e-6
m14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=28e-6
m15 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=433e-6
m16 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=13e-6
m17 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
m18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=237e-6
m19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=196e-6
m20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m21 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
m22 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
m23 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=237e-6
m24 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=467e-6
m25 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=467e-6
Capacitor1 outFirstStage out 10e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_80_9

** Expected Performance Values: 
** Gain: 110 dB
** Power consumption: 14.9991 mW
** Area: 12666 (mu_m)^2
** Transit frequency: 8.05401 MHz
** Transit frequency with error factor: 8.05366 MHz
** Slew rate: 30.3397 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** VoutMax: 4.25 V
** VoutMin: 1.17001 V
** VcmMax: 5.17001 V
** VcmMin: 1.96001 V


** Expected Currents: 
** NormalTransistorPmos: -9.93899e+06 muA
** NormalTransistorPmos: -1.68999e+07 muA
** NormalTransistorPmos: -5.37349e+07 muA
** NormalTransistorPmos: -3.07259e+08 muA
** NormalTransistorPmos: -4.7348e+08 muA
** NormalTransistorPmos: -3.07259e+08 muA
** NormalTransistorPmos: -4.7348e+08 muA
** NormalTransistorNmos: 3.0726e+08 muA
** NormalTransistorNmos: 3.07259e+08 muA
** NormalTransistorNmos: 3.0726e+08 muA
** NormalTransistorNmos: 3.07259e+08 muA
** NormalTransistorNmos: 3.3244e+08 muA
** DiodeTransistorNmos: 3.32439e+08 muA
** NormalTransistorNmos: 1.66221e+08 muA
** NormalTransistorNmos: 1.66221e+08 muA
** NormalTransistorNmos: 1.95237e+09 muA
** DiodeTransistorNmos: 1.95237e+09 muA
** NormalTransistorPmos: -1.95236e+09 muA
** DiodeTransistorNmos: 9.93801e+06 muA
** NormalTransistorNmos: 9.93701e+06 muA
** DiodeTransistorNmos: 1.68991e+07 muA
** NormalTransistorNmos: 1.68981e+07 muA
** DiodeTransistorNmos: 5.37341e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.31201  V
** outInputVoltageBiasXXnXX2: 1.57701  V
** outSourceVoltageBiasXXnXX1: 0.656001  V
** outSourceVoltageBiasXXnXX2: 0.790001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX3: 0.910001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.350001  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 4.23001  V
** sourceGCC2: 4.23001  V
** sourceTransconductance: 1.44401  V
** inner: 0.655001  V
** inner: 0.784001  V


.END