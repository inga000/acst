.suckt  two_stage_single_output_op_amp_9_12 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m3 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m4 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m5 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos
m6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c2 out sourceNmos 
m10 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m11 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m12 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m13 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
m14 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m16 ibias ibias sourceNmos sourceNmos nmos
m17 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m18 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_9_12

