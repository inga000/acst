** Name: two_stage_single_output_op_amp_110_3

.MACRO two_stage_single_output_op_amp_110_3 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=35e-6
m2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=101e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=101e-6
m4 ibias ibias outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos4 L=9e-6 W=49e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=32e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=121e-6
m7 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=9e-6 W=9e-6
m8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=5e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=181e-6
m10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=8e-6 W=101e-6
m11 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
m12 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=34e-6
m13 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=101e-6
m14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=9e-6 W=600e-6
m15 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=9e-6 W=59e-6
m16 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=4e-6
m17 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=121e-6
m18 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=4e-6
m19 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=98e-6
m20 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=98e-6
m21 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=9e-6 W=203e-6
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=32e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 7.30001e-12
.EOM two_stage_single_output_op_amp_110_3

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 2.30201 mW
** Area: 14988 (mu_m)^2
** Transit frequency: 2.81101 MHz
** Transit frequency with error factor: 2.8111 MHz
** Slew rate: 8.35538 V/mu_s
** Phase margin: 60.1606°
** CMRR: 127 dB
** VoutMax: 3.25 V
** VoutMin: 0.300001 V
** VcmMax: 3.04001 V
** VcmMin: 1.55001 V


** Expected Currents: 
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 6.54111e+07 muA
** NormalTransistorPmos: -6.67379e+07 muA
** NormalTransistorPmos: -2.40469e+07 muA
** NormalTransistorPmos: -2.40469e+07 muA
** DiodeTransistorNmos: 2.40461e+07 muA
** NormalTransistorNmos: 2.40461e+07 muA
** NormalTransistorNmos: 2.40461e+07 muA
** DiodeTransistorNmos: 2.40461e+07 muA
** NormalTransistorPmos: -1.13508e+08 muA
** DiodeTransistorPmos: -1.13509e+08 muA
** NormalTransistorPmos: -2.40479e+07 muA
** NormalTransistorPmos: -2.40479e+07 muA
** NormalTransistorNmos: 2.29627e+08 muA
** NormalTransistorPmos: -2.29626e+08 muA
** NormalTransistorPmos: -2.29625e+08 muA
** DiodeTransistorNmos: 6.67371e+07 muA
** DiodeTransistorPmos: -3.04759e+07 muA
** NormalTransistorPmos: -3.04769e+07 muA
** DiodeTransistorPmos: -6.54119e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.79901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outInputVoltageBiasXXpXX1: 3.41201  V
** outSourceVoltageBiasXXpXX1: 4.20601  V
** outSourceVoltageBiasXXpXX3: 3.68501  V
** outVoltageBiasXXpXX2: 1.39401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.43301  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 2.96701  V
** sourceGCC2: 2.95801  V
** innerStageBias: 3.80001  V
** inner: 4.20601  V


.END