.suckt  two_stage_fully_differential_op_amp_13_1 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_Load_2 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_3 outFeedback outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_4 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_5 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackStage_Transconductor_6 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_7 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_8 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FeedbackStage_Transconductor_9 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FirstStage_Load_10 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_11 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_StageBias_12 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Transconductor_13 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_FullyDifferential_FirstStage_Transconductor_14 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_Transconductor_15 out1 out1FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_16 out1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_Transconductor_17 out2 out2FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_StageBias_18 out2 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_19 ibias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_20 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_13_1

