.suckt  complementary_op_amp19 ibias in1 in2 out sourceNmos sourcePmos
m_Complementary_MainBias_1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_2 FirstStageYinnerOutputLoadNmos FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m_Complementary_FirstStage_Load_3 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerOutputLoadNmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_4 out FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m_Complementary_FirstStage_Load_5 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerOutputLoadNmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_6 FirstStageYinnerOutputLoadNmos FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m_Complementary_FirstStage_Load_7 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerOutputLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_8 out FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m_Complementary_FirstStage_Load_9 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerOutputLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_10 FirstStageYsourceTransconductanceNmos outInputVoltageBiasXXnXX1 FirstStageYinnerStageBiasNmos FirstStageYinnerStageBiasNmos nmos
m_Complementary_FirstStage_StageBias_11 FirstStageYinnerStageBiasNmos outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_12 FirstStageYsourceTransconductancePmos ibias FirstStageYinnerStageBiasPmos FirstStageYinnerStageBiasPmos pmos
m_Complementary_FirstStage_StageBias_13 FirstStageYinnerStageBiasPmos outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Transconductor_14 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_15 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_16 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m_Complementary_FirstStage_Transconductor_17 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c_Complementary_Load_Capacitor_1 out sourceNmos 
m_Complementary_MainBias_18 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_Complementary_MainBias_19 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_MainBias_20 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_Complementary_MainBias_21 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end complementary_op_amp19

