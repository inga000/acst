** Name: two_stage_single_output_op_amp_68_1

.MACRO two_stage_single_output_op_amp_68_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=33e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=47e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=7e-6 W=14e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=14e-6
mMainBias5 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=12e-6
mMainBias6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=8e-6 W=39e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=205e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=9e-6 W=42e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=119e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=119e-6
mMainBias11 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=82e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=253e-6
mFoldedCascodeFirstStageLoad13 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=9e-6 W=42e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=15e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=7e-6 W=14e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=15e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=15e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=8e-6 W=205e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=39e-6
mSecondStage1StageBias20 out inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=461e-6
mFoldedCascodeFirstStageLoad21 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=14e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_68_1

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 3.70201 mW
** Area: 12345 (mu_m)^2
** Transit frequency: 3.34701 MHz
** Transit frequency with error factor: 3.34713 MHz
** Slew rate: 3.70858 V/mu_s
** Phase margin: 61.3065°
** CMRR: 139 dB
** VoutMax: 4.51001 V
** VoutMin: 0.530001 V
** VcmMax: 3.31001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.17801e+06 muA
** NormalTransistorNmos: 1.74761e+07 muA
** NormalTransistorNmos: 1.67601e+07 muA
** NormalTransistorNmos: 2.51841e+07 muA
** NormalTransistorNmos: 1.67601e+07 muA
** NormalTransistorNmos: 2.51841e+07 muA
** DiodeTransistorPmos: -1.67609e+07 muA
** NormalTransistorPmos: -1.67619e+07 muA
** NormalTransistorPmos: -1.67609e+07 muA
** DiodeTransistorPmos: -1.67619e+07 muA
** NormalTransistorPmos: -1.68509e+07 muA
** DiodeTransistorPmos: -1.68519e+07 muA
** NormalTransistorPmos: -8.42499e+06 muA
** NormalTransistorPmos: -8.42499e+06 muA
** NormalTransistorNmos: 6.59319e+08 muA
** NormalTransistorPmos: -6.59318e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.17899e+06 muA
** NormalTransistorPmos: -3.17999e+06 muA
** DiodeTransistorPmos: -1.74769e+07 muA


** Expected Voltages: 
** ibias: 1.13901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.94401  V
** out: 2.5  V
** outFirstStage: 0.934001  V
** outInputVoltageBiasXXpXX1: 3.48801  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.24401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 3.74601  V
** innerTransistorStack2Load2: 3.74801  V
** out1: 2.92401  V
** sourceGCC1: 0.527001  V
** sourceGCC2: 0.527001  V
** sourceTransconductance: 3.24101  V
** inner: 4.24301  V


.END