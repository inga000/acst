** Name: two_stage_single_output_op_amp_9_9

.MACRO two_stage_single_output_op_amp_9_9 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=25e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=7e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=125e-6
m4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=51e-6
m5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
m6 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=125e-6
m7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=21e-6
m8 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=45e-6
m9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=21e-6
m10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=9e-6 W=106e-6
m11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
m12 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=212e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=538e-6
m14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=42e-6
m15 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 5.30001e-12
.EOM two_stage_single_output_op_amp_9_9

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 7.44801 mW
** Area: 5452 (mu_m)^2
** Transit frequency: 8.19701 MHz
** Transit frequency with error factor: 8.19127 MHz
** Slew rate: 7.9339 V/mu_s
** Phase margin: 60.1606°
** CMRR: 102 dB
** negPSRR: 102 dB
** posPSRR: 94 dB
** VoutMax: 4.25 V
** VoutMin: 1.63001 V
** VcmMax: 4.32001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorNmos: 1.80441e+07 muA
** NormalTransistorPmos: -7.39679e+07 muA
** NormalTransistorPmos: -2.10949e+07 muA
** NormalTransistorPmos: -2.10949e+07 muA
** DiodeTransistorPmos: -2.10949e+07 muA
** NormalTransistorNmos: 4.21871e+07 muA
** NormalTransistorNmos: 2.10941e+07 muA
** NormalTransistorNmos: 2.10941e+07 muA
** NormalTransistorNmos: 1.34536e+09 muA
** DiodeTransistorNmos: 1.34536e+09 muA
** NormalTransistorPmos: -1.34535e+09 muA
** DiodeTransistorNmos: 7.39671e+07 muA
** NormalTransistorNmos: 7.39671e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.80449e+07 muA


** Expected Voltages: 
** ibias: 0.611001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.04001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 1.02001  V
** outVoltageBiasXXpXX0: 4.23801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.28601  V
** out1: 3.34901  V
** sourceTransconductance: 1.94101  V
** inner: 1.02001  V


.END