.suckt  symmetrical_op_amp54 ibias in1 in2 out sourceNmos sourcePmos
mSymmetricalFirstStageLoad1 outFirstStage outFirstStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageLoad2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageStageBias3 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mSymmetricalFirstStageStageBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mSymmetricalFirstStageTransconductor5 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSymmetricalFirstStageTransconductor6 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias8 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos
mSecondStage1StageBias9 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias10 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias11 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor12 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mMainBias13 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mMainBias14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end symmetrical_op_amp54

