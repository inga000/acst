.suckt  two_stage_fully_differential_op_amp_6_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_3 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_Load_5 outFeedback outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_6 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_8 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackStage_Transconductor_10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FeedbackStage_Transconductor_13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FirstStage_Load_14 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m_FullyDifferential_FirstStage_Load_15 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_16 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m_FullyDifferential_FirstStage_Load_17 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_18 out1FirstStage ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_19 out2FirstStage ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_StageBias_20 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Transconductor_21 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_FullyDifferential_FirstStage_Transconductor_22 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_Transconductor_23 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m_FullyDifferential_SecondStage1_Transconductor_24 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_25 out1 outVoltageBiasXXpXX1 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m_FullyDifferential_SecondStage1_StageBias_26 SecondStage1YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_Transconductor_27 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m_FullyDifferential_SecondStage2_Transconductor_28 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_StageBias_29 out2 outVoltageBiasXXpXX1 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m_FullyDifferential_SecondStage2_StageBias_30 SecondStage2YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_31 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_32 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_33 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_34 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_6_4

