** Name: two_stage_single_output_op_amp_39_7

.MACRO two_stage_single_output_op_amp_39_7 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=22e-6
m3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=41e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=41e-6
m5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=36e-6
m6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=26e-6
m7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=7e-6
m8 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=8e-6 W=10e-6
m9 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=546e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=7e-6
m11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=16e-6
m12 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=41e-6
m13 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=252e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=292e-6
m15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=41e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_39_7

** Expected Performance Values: 
** Gain: 84 dB
** Power consumption: 2.76101 mW
** Area: 6585 (mu_m)^2
** Transit frequency: 2.70801 MHz
** Transit frequency with error factor: 2.70469 MHz
** Slew rate: 4.40966 V/mu_s
** Phase margin: 60.7336°
** CMRR: 102 dB
** negPSRR: 94 dB
** posPSRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 0.160001 V
** VcmMax: 3.91001 V
** VcmMin: 1.67001 V


** Expected Currents: 
** NormalTransistorNmos: 1.21701e+07 muA
** NormalTransistorPmos: -8.65719e+07 muA
** DiodeTransistorPmos: -9.95299e+06 muA
** NormalTransistorPmos: -9.95199e+06 muA
** NormalTransistorPmos: -9.95299e+06 muA
** DiodeTransistorPmos: -9.95199e+06 muA
** NormalTransistorNmos: 1.99031e+07 muA
** NormalTransistorNmos: 1.99021e+07 muA
** NormalTransistorNmos: 9.95201e+06 muA
** NormalTransistorNmos: 9.95201e+06 muA
** NormalTransistorNmos: 4.23542e+08 muA
** NormalTransistorPmos: -4.23541e+08 muA
** DiodeTransistorNmos: 8.65711e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.21709e+07 muA


** Expected Voltages: 
** ibias: 0.570001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.01201  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 4.07101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.27201  V
** innerStageBias: 0.172001  V
** innerTransistorStack1Load1: 4.27201  V
** out1: 3.50701  V
** sourceTransconductance: 1.83501  V


.END