** Name: two_stage_single_output_op_amp_187_9

.MACRO two_stage_single_output_op_amp_187_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=6e-6
m2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=1e-6 W=25e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=407e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=54e-6
m5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
m6 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=43e-6
m7 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=407e-6
m8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=7e-6 W=8e-6
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=16e-6
m10 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=30e-6
m11 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=9e-6
m12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=16e-6
m13 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=29e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
m15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=104e-6
m16 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=467e-6
m17 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=502e-6
m18 outFirstStage ibias sourcePmos sourcePmos pmos4 L=2e-6 W=358e-6
m19 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=358e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.90001e-12
.EOM two_stage_single_output_op_amp_187_9

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 10.1161 mW
** Area: 6116 (mu_m)^2
** Transit frequency: 6.47301 MHz
** Transit frequency with error factor: 6.45906 MHz
** Slew rate: 6.10051 V/mu_s
** Phase margin: 60.1606°
** CMRR: 88 dB
** VoutMax: 4.25 V
** VoutMin: 1.03001 V
** VcmMax: 5.24001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorPmos: -2.46329e+07 muA
** NormalTransistorPmos: -1.10612e+08 muA
** NormalTransistorNmos: 5.39761e+07 muA
** NormalTransistorNmos: 5.39751e+07 muA
** DiodeTransistorNmos: 5.39761e+07 muA
** NormalTransistorPmos: -8.44509e+07 muA
** NormalTransistorPmos: -8.44509e+07 muA
** NormalTransistorNmos: 6.09491e+07 muA
** NormalTransistorNmos: 6.09481e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 1.69901e+09 muA
** DiodeTransistorNmos: 1.69901e+09 muA
** NormalTransistorPmos: -1.699e+09 muA
** DiodeTransistorNmos: 2.46321e+07 muA
** NormalTransistorNmos: 2.46331e+07 muA
** DiodeTransistorNmos: 1.10613e+08 muA
** DiodeTransistorNmos: 1.10612e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.43601  V
** inputVoltageBiasXXnXX2: 1.19301  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.718001  V
** outSourceVoltageBiasXXnXX2: 0.560001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.940001  V
** innerStageBias: 0.630001  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 0.719001  V


.END