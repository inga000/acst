** Name: two_stage_single_output_op_amp_81_7

.MACRO two_stage_single_output_op_amp_81_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=9e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=39e-6
m5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m7 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=331e-6
m8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=3e-6 W=39e-6
m9 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
m10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=39e-6
m11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=24e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=24e-6
m13 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=25e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=197e-6
m15 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=102e-6
m16 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=447e-6
m17 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=54e-6
m18 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=102e-6
m19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
m20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_81_7

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 13.2701 mW
** Area: 2270 (mu_m)^2
** Transit frequency: 11.0591 MHz
** Transit frequency with error factor: 11.0587 MHz
** Slew rate: 9.12736 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 0.380001 V
** VcmMax: 5.17001 V
** VcmMin: 1.5 V


** Expected Currents: 
** NormalTransistorPmos: -4.47858e+08 muA
** NormalTransistorPmos: -5.41759e+07 muA
** NormalTransistorPmos: -4.14249e+07 muA
** NormalTransistorPmos: -6.59019e+07 muA
** NormalTransistorPmos: -4.14249e+07 muA
** NormalTransistorPmos: -6.59019e+07 muA
** DiodeTransistorNmos: 4.14241e+07 muA
** NormalTransistorNmos: 4.14231e+07 muA
** NormalTransistorNmos: 4.14241e+07 muA
** DiodeTransistorNmos: 4.14231e+07 muA
** NormalTransistorNmos: 4.89511e+07 muA
** NormalTransistorNmos: 4.89501e+07 muA
** NormalTransistorNmos: 2.44761e+07 muA
** NormalTransistorNmos: 2.44761e+07 muA
** NormalTransistorNmos: 2.00023e+09 muA
** NormalTransistorPmos: -2.00022e+09 muA
** DiodeTransistorNmos: 4.47859e+08 muA
** DiodeTransistorNmos: 5.41751e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.13601  V
** outVoltageBiasXXnXX2: 0.784001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.563001  V
** innerStageBias: 0.579001  V
** innerTransistorStack1Load2: 0.563001  V
** out1: 1.16201  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.93901  V


.END