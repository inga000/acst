.suckt  two_stage_single_output_op_amp_192_10 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_4 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_6 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m_SingleOutput_FirstStage_Load_7 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_8 FirstStageYout1 ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_9 outFirstStage ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_StageBias_10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_SingleOutput_FirstStage_StageBias_11 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Transconductor_12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_SingleOutput_FirstStage_Transconductor_13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_StageBias_14 out inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_Transconductor_15 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m_SingleOutput_SecondStage1_Transconductor_16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_17 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_SingleOutput_MainBias_18 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_19 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_20 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_21 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_22 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_192_10

