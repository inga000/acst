** Name: two_stage_single_output_op_amp_24_2

.MACRO two_stage_single_output_op_amp_24_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=12e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=22e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=18e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=221e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=439e-6
m6 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=7e-6 W=411e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=128e-6
m8 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=49e-6
m9 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=128e-6
m10 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=108e-6
m11 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=108e-6
m12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=201e-6
m13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=31e-6
m14 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=340e-6
m15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=116e-6
m16 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=34e-6
m17 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=116e-6
m18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=439e-6
m19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=221e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10.6001e-12
.EOM two_stage_single_output_op_amp_24_2

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 1.86501 mW
** Area: 13907 (mu_m)^2
** Transit frequency: 2.91001 MHz
** Transit frequency with error factor: 2.90606 MHz
** Slew rate: 6.22781 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** negPSRR: 97 dB
** posPSRR: 111 dB
** VoutMax: 4.69001 V
** VoutMin: 0.350001 V
** VcmMax: 3.09001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.21291e+07 muA
** NormalTransistorPmos: -1.91549e+07 muA
** NormalTransistorPmos: -1.74649e+07 muA
** NormalTransistorNmos: 4.13331e+07 muA
** NormalTransistorNmos: 4.13321e+07 muA
** NormalTransistorNmos: 4.13331e+07 muA
** NormalTransistorNmos: 4.13321e+07 muA
** NormalTransistorPmos: -8.26689e+07 muA
** DiodeTransistorPmos: -8.26699e+07 muA
** NormalTransistorPmos: -4.13339e+07 muA
** NormalTransistorPmos: -4.13339e+07 muA
** NormalTransistorNmos: 1.91553e+08 muA
** NormalTransistorNmos: 1.91552e+08 muA
** NormalTransistorPmos: -1.91552e+08 muA
** DiodeTransistorNmos: 1.91541e+07 muA
** DiodeTransistorNmos: 1.74641e+07 muA
** DiodeTransistorPmos: -4.21299e+07 muA
** NormalTransistorPmos: -4.21299e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.751001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.51601  V
** outSourceVoltageBiasXXpXX1: 4.25801  V
** outVoltageBiasXXnXX0: 0.631001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.182001  V
** innerTransistorStack2Load1: 0.182001  V
** sourceTransconductance: 3.48601  V
** innerTransconductance: 0.150001  V
** inner: 4.25801  V


.END