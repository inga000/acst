** Name: symmetrical_op_amp81

.MACRO symmetrical_op_amp81 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=19e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=600e-6
mSecondStage1StageBias4 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=7e-6
mSymmetricalFirstStageLoad5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=193e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=9e-6
mSymmetricalFirstStageLoad7 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=193e-6
mSymmetricalFirstStageStageBias8 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=600e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=78e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias10 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=78e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=19e-6
mMainBias12 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=19e-6
mSymmetricalFirstStageTransconductor13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=58e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias14 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=1e-6 W=68e-6
mMainBias15 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=18e-6
mSecondStage1StageBias16 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=68e-6
mSymmetricalFirstStageTransconductor17 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=58e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=183e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor19 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=183e-6
mMainBias20 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=9e-6 W=76e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor21 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=7e-6 W=209e-6
mSecondStage1Transconductor22 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=7e-6 W=209e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp81

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 3.60701 mW
** Area: 14647 (mu_m)^2
** Transit frequency: 4.64901 MHz
** Transit frequency with error factor: 4.64876 MHz
** Slew rate: 14.9439 V/mu_s
** Phase margin: 70.4739°
** CMRR: 135 dB
** negPSRR: 41 dB
** posPSRR: 35 dB
** VoutMax: 4.26001 V
** VoutMin: 0.310001 V
** VcmMax: 4.63001 V
** VcmMin: 1.73001 V


** Expected Currents: 
** NormalTransistorNmos: 9.44901e+06 muA
** NormalTransistorNmos: 1.00401e+07 muA
** NormalTransistorPmos: -8.12279e+07 muA
** DiodeTransistorPmos: -1.55507e+08 muA
** DiodeTransistorPmos: -1.55507e+08 muA
** NormalTransistorNmos: 3.11014e+08 muA
** DiodeTransistorNmos: 3.11013e+08 muA
** NormalTransistorNmos: 1.55508e+08 muA
** NormalTransistorNmos: 1.55508e+08 muA
** NormalTransistorNmos: 1.49865e+08 muA
** NormalTransistorNmos: 1.49864e+08 muA
** NormalTransistorPmos: -1.49864e+08 muA
** NormalTransistorPmos: -1.49863e+08 muA
** NormalTransistorNmos: 1.49865e+08 muA
** NormalTransistorNmos: 1.49864e+08 muA
** NormalTransistorPmos: -1.49864e+08 muA
** NormalTransistorPmos: -1.49863e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 8.12271e+07 muA
** DiodeTransistorPmos: -9.44999e+06 muA
** DiodeTransistorPmos: -1.00409e+07 muA


** Expected Voltages: 
** ibias: 1.22401  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.716001  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 4.22301  V
** innerComplementarySecondStage: 0.555001  V
** inputVoltageBiasXXpXX0: 3.70601  V
** out: 2.5  V
** outFirstStage: 4.22301  V
** outSourceVoltageBiasXXnXX1: 0.613001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.59001  V
** innerStageBias: 0.150001  V
** innerTransconductance: 4.77801  V
** inner: 0.150001  V
** inner: 4.77801  V
** inner: 0.610001  V


.END