.suckt  two_stage_single_output_op_amp_175_10 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mMainBias2 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad5 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos
mSimpleFirstStageLoad6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad7 FirstStageYout1 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad8 outFirstStage ibias sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias13 out ibias sourceNmos sourceNmos nmos
mSecondStage1Transconductor14 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor15 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
mMainBias16 ibias ibias sourceNmos sourceNmos nmos
mSecondStage1StageBias17 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mMainBias18 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_175_10

