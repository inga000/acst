.suckt  symmetrical_op_amp37 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mMainBias2 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
mMainBias3 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad4 outFirstStage outFirstStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageLoad5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
mSymmetricalFirstStageStageBias7 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos
mSymmetricalFirstStageTransconductor8 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1Transconductor10 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mSecondStage1Transconductor11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias12 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mSecondStage1StageBias13 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias14 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias15 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mMainBias18 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
mSecondStage1StageBias19 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
mMainBias20 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
mMainBias21 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp37

