** Name: two_stage_single_output_op_amp_64_2

.MACRO two_stage_single_output_op_amp_64_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=9e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
m3 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=10e-6
m4 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=18e-6
m6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=11e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=203e-6
m8 FirstStageYinnerOutputLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=202e-6
m9 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=344e-6
m10 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=344e-6
m11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=496e-6
m12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=600e-6
m13 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=202e-6
m14 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=16e-6
m15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=151e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=151e-6
m18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=203e-6
m19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m20 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=8e-6
m21 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=576e-6
m22 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=10e-6
m23 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=48e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 18.4001e-12
.EOM two_stage_single_output_op_amp_64_2

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 3.63101 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 2.85401 MHz
** Transit frequency with error factor: 2.85435 MHz
** Slew rate: 5.4011 V/mu_s
** Phase margin: 60.1606°
** CMRR: 118 dB
** VoutMax: 4.75 V
** VoutMin: 0.350001 V
** VcmMax: 3.05001 V
** VcmMin: -0.389999 V


** Expected Currents: 
** NormalTransistorNmos: 7.86001e+06 muA
** NormalTransistorPmos: -2.66239e+07 muA
** NormalTransistorPmos: -4.42399e+06 muA
** NormalTransistorNmos: 9.98871e+07 muA
** NormalTransistorNmos: 1.71237e+08 muA
** NormalTransistorNmos: 9.98831e+07 muA
** NormalTransistorNmos: 1.71231e+08 muA
** DiodeTransistorPmos: -9.98859e+07 muA
** DiodeTransistorPmos: -9.98849e+07 muA
** NormalTransistorPmos: -9.98839e+07 muA
** NormalTransistorPmos: -9.98849e+07 muA
** NormalTransistorPmos: -1.42696e+08 muA
** DiodeTransistorPmos: -1.42697e+08 muA
** NormalTransistorPmos: -7.13479e+07 muA
** NormalTransistorPmos: -7.13479e+07 muA
** NormalTransistorNmos: 3.24909e+08 muA
** NormalTransistorNmos: 3.24908e+08 muA
** NormalTransistorPmos: -3.24908e+08 muA
** DiodeTransistorNmos: 2.66231e+07 muA
** DiodeTransistorNmos: 4.42301e+06 muA
** DiodeTransistorPmos: -7.86099e+06 muA
** NormalTransistorPmos: -7.86199e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.576001  V
** out: 2.5  V
** outFirstStage: 0.558001  V
** outInputVoltageBiasXXpXX1: 3.47401  V
** outSourceVoltageBiasXXpXX1: 4.23701  V
** outVoltageBiasXXnXX1: 0.963001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 2.43701  V
** innerTransistorStack1Load2: 3.75101  V
** innerTransistorStack2Load2: 3.74501  V
** sourceGCC1: 0.371001  V
** sourceGCC2: 0.371001  V
** sourceTransconductance: 3.49301  V
** innerTransconductance: 0.362001  V
** inner: 4.23701  V


.END