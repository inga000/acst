** Name: two_stage_single_output_op_amp_90_1

.MACRO two_stage_single_output_op_amp_90_1 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=148e-6
mTelescopicFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=148e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=6e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=34e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=148e-6
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=279e-6
mTelescopicFirstStageLoad8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=9e-6 W=148e-6
mMainBias9 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=4e-6 W=24e-6
mTelescopicFirstStageLoad10 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=129e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=9e-6 W=332e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=9e-6 W=332e-6
mMainBias13 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
mSecondStage1StageBias14 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=523e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=129e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=98e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 15.2001e-12
.EOM two_stage_single_output_op_amp_90_1

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 3.27601 mW
** Area: 14988 (mu_m)^2
** Transit frequency: 2.99001 MHz
** Transit frequency with error factor: 2.99049 MHz
** Slew rate: 6.52849 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.66001 V
** VoutMin: 0.300001 V
** VcmMax: 3.88001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorNmos: 3.72071e+07 muA
** NormalTransistorPmos: -9.16999e+06 muA
** NormalTransistorPmos: -3.13219e+07 muA
** NormalTransistorPmos: -3.13219e+07 muA
** DiodeTransistorNmos: 3.13211e+07 muA
** NormalTransistorNmos: 3.13211e+07 muA
** NormalTransistorNmos: 3.13211e+07 muA
** DiodeTransistorNmos: 3.13211e+07 muA
** NormalTransistorPmos: -9.98529e+07 muA
** NormalTransistorPmos: -3.13229e+07 muA
** NormalTransistorPmos: -3.13229e+07 muA
** NormalTransistorNmos: 5.26131e+08 muA
** NormalTransistorPmos: -5.2613e+08 muA
** DiodeTransistorNmos: 9.16901e+06 muA
** DiodeTransistorPmos: -3.72079e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.10001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.675001  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outVoltageBiasXXpXX1: 2.22001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.28101  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 3.01601  V
** sourceGCC2: 3.01601  V


.END