** Name: two_stage_single_output_op_amp_47_10

.MACRO two_stage_single_output_op_amp_47_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=41e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=81e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=86e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=86e-6
mMainBias8 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=79e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=598e-6
mFoldedCascodeFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=81e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=77e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=199e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=199e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=228e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=228e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=600e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=519e-6
mMainBias18 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=123e-6
mSecondStage1Transconductor19 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=77e-6
mMainBias21 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=406e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 16.6001e-12
.EOM two_stage_single_output_op_amp_47_10

** Expected Performance Values: 
** Gain: 131 dB
** Power consumption: 10.6941 mW
** Area: 8659 (mu_m)^2
** Transit frequency: 7.43501 MHz
** Transit frequency with error factor: 7.43461 MHz
** Slew rate: 7.48252 V/mu_s
** Phase margin: 60.1606°
** CMRR: 140 dB
** VoutMax: 4.25 V
** VoutMin: 0.170001 V
** VcmMax: 4.01001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorNmos: 1.82761e+08 muA
** NormalTransistorPmos: -1.00318e+08 muA
** NormalTransistorPmos: -3.00249e+07 muA
** NormalTransistorNmos: 1.24493e+08 muA
** NormalTransistorNmos: 1.9862e+08 muA
** NormalTransistorNmos: 1.24493e+08 muA
** NormalTransistorNmos: 1.9862e+08 muA
** NormalTransistorPmos: -1.24492e+08 muA
** NormalTransistorPmos: -1.24493e+08 muA
** NormalTransistorPmos: -1.24492e+08 muA
** NormalTransistorPmos: -1.24493e+08 muA
** NormalTransistorPmos: -1.48254e+08 muA
** NormalTransistorPmos: -7.41279e+07 muA
** NormalTransistorPmos: -7.41279e+07 muA
** NormalTransistorNmos: 1.40844e+09 muA
** NormalTransistorPmos: -1.40843e+09 muA
** NormalTransistorPmos: -1.40843e+09 muA
** DiodeTransistorNmos: 1.00319e+08 muA
** DiodeTransistorNmos: 3.00241e+07 muA
** DiodeTransistorPmos: -1.8276e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.20201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.571001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.04701  V
** outVoltageBiasXXnXX1: 1.00401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.24801  V
** innerTransistorStack1Load2: 4.55001  V
** innerTransistorStack2Load2: 4.55001  V
** sourceGCC1: 0.366001  V
** sourceGCC2: 0.366001  V
** sourceTransconductance: 3.25401  V
** innerTransconductance: 4.61101  V


.END