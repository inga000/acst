** Name: two_stage_single_output_op_amp_44_9

.MACRO two_stage_single_output_op_amp_44_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=4e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=5e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=433e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=57e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=121e-6
m6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
m7 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=433e-6
m8 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=4e-6
m9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=4e-6
m10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=93e-6
m11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=93e-6
m12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=94e-6
m14 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=439e-6
m15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=3e-6 W=94e-6
m16 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=131e-6
m17 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=27e-6
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=79e-6
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=79e-6
m20 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=7e-6 W=479e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_44_9

** Expected Performance Values: 
** Gain: 112 dB
** Power consumption: 5.60401 mW
** Area: 12961 (mu_m)^2
** Transit frequency: 4.79101 MHz
** Transit frequency with error factor: 4.79072 MHz
** Slew rate: 8.67692 V/mu_s
** Phase margin: 64.7443°
** CMRR: 127 dB
** VoutMax: 4.25 V
** VoutMin: 0.960001 V
** VcmMax: 3.97001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.08569e+07 muA
** NormalTransistorPmos: -3.61879e+07 muA
** NormalTransistorNmos: 3.92971e+07 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorNmos: 3.92971e+07 muA
** NormalTransistorNmos: 5.90441e+07 muA
** NormalTransistorPmos: -3.92979e+07 muA
** NormalTransistorPmos: -3.92979e+07 muA
** DiodeTransistorPmos: -3.92979e+07 muA
** NormalTransistorPmos: -3.94969e+07 muA
** NormalTransistorPmos: -1.97479e+07 muA
** NormalTransistorPmos: -1.97479e+07 muA
** NormalTransistorNmos: 9.35668e+08 muA
** DiodeTransistorNmos: 9.35667e+08 muA
** NormalTransistorPmos: -9.35667e+08 muA
** DiodeTransistorNmos: 1.08561e+07 muA
** NormalTransistorNmos: 1.08551e+07 muA
** DiodeTransistorNmos: 3.61871e+07 muA
** DiodeTransistorNmos: 3.61881e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.52401  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.36201  V
** outSourceVoltageBiasXXnXX1: 0.681001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.15001  V
** out1: 3.32201  V
** sourceGCC1: 0.526001  V
** sourceGCC2: 0.526001  V
** sourceTransconductance: 3.35301  V
** inner: 0.679001  V


.END