** Name: two_stage_single_output_op_amp_78_1

.MACRO two_stage_single_output_op_amp_78_1 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=86e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=64e-6
mMainBias3 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=50e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=116e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=5e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourceNmos sourceNmos nmos4 L=9e-6 W=86e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=7e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=116e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=50e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=137e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=64e-6
mMainBias14 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=85e-6
mMainBias15 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=102e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=31e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=551e-6
mFoldedCascodeFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=31e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_78_1

** Expected Performance Values: 
** Gain: 118 dB
** Power consumption: 3.16001 mW
** Area: 9575 (mu_m)^2
** Transit frequency: 3.90701 MHz
** Transit frequency with error factor: 3.90647 MHz
** Slew rate: 3.84691 V/mu_s
** Phase margin: 60.1606°
** CMRR: 139 dB
** VoutMax: 4.77001 V
** VoutMin: 0.520001 V
** VcmMax: 5.17001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 1.69211e+07 muA
** NormalTransistorNmos: 2.04011e+07 muA
** NormalTransistorPmos: -1.81999e+07 muA
** NormalTransistorPmos: -2.95799e+07 muA
** NormalTransistorPmos: -1.81999e+07 muA
** NormalTransistorPmos: -2.95799e+07 muA
** DiodeTransistorNmos: 1.81991e+07 muA
** DiodeTransistorNmos: 1.82001e+07 muA
** NormalTransistorNmos: 1.81991e+07 muA
** NormalTransistorNmos: 1.82001e+07 muA
** NormalTransistorNmos: 2.27581e+07 muA
** DiodeTransistorNmos: 2.27591e+07 muA
** NormalTransistorNmos: 1.13791e+07 muA
** NormalTransistorNmos: 1.13791e+07 muA
** NormalTransistorNmos: 5.25459e+08 muA
** NormalTransistorPmos: -5.25458e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.69219e+07 muA
** DiodeTransistorPmos: -2.04019e+07 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.929001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.20401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.555001  V
** innerTransistorStack2Load2: 0.555001  V
** out1: 1.13401  V
** sourceGCC1: 4.56301  V
** sourceGCC2: 4.56301  V
** sourceTransconductance: 1.89901  V
** inner: 0.556001  V


.END