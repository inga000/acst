.suckt  two_stage_single_output_op_amp_1_7 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad3 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias7 out outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mSecondStage1Transconductor8 out outFirstStage sourcePmos sourcePmos pmos
mMainBias9 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias10 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_1_7

