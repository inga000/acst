** Name: two_stage_single_output_op_amp_31_9

.MACRO two_stage_single_output_op_amp_31_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=7e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=198e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=113e-6
mMainBias6 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mSimpleFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=93e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=54e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=48e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=10e-6
mMainBias11 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=198e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=54e-6
mSimpleFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=113e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=533e-6
mSimpleFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=68e-6
mMainBias17 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=77e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.30001e-12
.EOM two_stage_single_output_op_amp_31_9

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 10.0341 mW
** Area: 4155 (mu_m)^2
** Transit frequency: 8.73301 MHz
** Transit frequency with error factor: 8.72629 MHz
** Slew rate: 10.9776 V/mu_s
** Phase margin: 60.1606°
** CMRR: 102 dB
** negPSRR: 95 dB
** posPSRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 1.54001 V
** VcmMax: 4.42001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 1.18261e+07 muA
** NormalTransistorPmos: -8.95e+07 muA
** NormalTransistorPmos: -4.57389e+07 muA
** NormalTransistorPmos: -4.57389e+07 muA
** DiodeTransistorPmos: -4.57389e+07 muA
** NormalTransistorNmos: 9.14751e+07 muA
** NormalTransistorNmos: 9.14741e+07 muA
** NormalTransistorNmos: 4.57381e+07 muA
** NormalTransistorNmos: 4.57381e+07 muA
** NormalTransistorNmos: 1.80393e+09 muA
** DiodeTransistorNmos: 1.80393e+09 muA
** NormalTransistorPmos: -1.80392e+09 muA
** DiodeTransistorNmos: 8.94991e+07 muA
** NormalTransistorNmos: 8.94991e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.18269e+07 muA


** Expected Voltages: 
** ibias: 1.14601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.07401  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.94201  V
** outSourceVoltageBiasXXnXX1: 0.971001  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.28601  V
** innerStageBias: 0.528001  V
** out1: 3.44901  V
** sourceTransconductance: 1.89401  V
** inner: 0.971001  V


.END