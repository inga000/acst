** Name: two_stage_single_output_op_amp_48_7

.MACRO two_stage_single_output_op_amp_48_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=10e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=64e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=264e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=264e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=9e-6 W=83e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=99e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=99e-6
mSecondStage1StageBias9 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad10 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=9e-6 W=83e-6
mFoldedCascodeFirstStageLoad11 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=264e-6
mFoldedCascodeFirstStageTransconductor12 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=74e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=74e-6
mFoldedCascodeFirstStageStageBias14 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=600e-6
mSecondStage1Transconductor15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=244e-6
mFoldedCascodeFirstStageLoad16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=264e-6
mMainBias17 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=196e-6
mMainBias18 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=481e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 20.4001e-12
.EOM two_stage_single_output_op_amp_48_7

** Expected Performance Values: 
** Gain: 114 dB
** Power consumption: 8.61301 mW
** Area: 9310 (mu_m)^2
** Transit frequency: 3.48201 MHz
** Transit frequency with error factor: 3.48201 MHz
** Slew rate: 5.48927 V/mu_s
** Phase margin: 60.1606°
** CMRR: 133 dB
** VoutMax: 4.48001 V
** VoutMin: 0.150001 V
** VcmMax: 3.86001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -4.93559e+07 muA
** NormalTransistorPmos: -1.21897e+08 muA
** NormalTransistorNmos: 1.12517e+08 muA
** NormalTransistorNmos: 1.88559e+08 muA
** NormalTransistorNmos: 1.12517e+08 muA
** NormalTransistorNmos: 1.88559e+08 muA
** DiodeTransistorPmos: -1.12516e+08 muA
** NormalTransistorPmos: -1.12517e+08 muA
** NormalTransistorPmos: -1.12516e+08 muA
** DiodeTransistorPmos: -1.12517e+08 muA
** NormalTransistorPmos: -1.5208e+08 muA
** NormalTransistorPmos: -7.60409e+07 muA
** NormalTransistorPmos: -7.60409e+07 muA
** NormalTransistorNmos: 1.15432e+09 muA
** NormalTransistorPmos: -1.15431e+09 muA
** DiodeTransistorNmos: 4.93551e+07 muA
** DiodeTransistorNmos: 1.21898e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.91901  V
** outVoltageBiasXXnXX1: 1.13301  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.28101  V
** innerTransistorStack1Load2: 4.28001  V
** out1: 3.56201  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.40201  V


.END