.suckt  two_stage_fully_differential_op_amp_67_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m2 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m3 outVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m4 inputVoltageBiasXXnXX4 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m5 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m6 outFeedback outFeedback sourcePmos sourcePmos pmos
m7 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m8 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m9 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 out1FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m14 out2FirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m15 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m16 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m17 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m18 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m19 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m20 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m21 out1 outVoltageBiasXXnXX3 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m22 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m23 out1 ibias SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m24 SecondStage1YinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m25 out2 outVoltageBiasXXnXX3 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m26 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m27 out2 ibias SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m28 SecondStage2YinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m29 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m30 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m31 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos
m32 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m33 inputVoltageBiasXXnXX4 inputVoltageBiasXXnXX4 sourceNmos sourceNmos nmos
m34 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m35 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_67_4

