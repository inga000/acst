** Name: symmetrical_op_amp83

.MACRO symmetrical_op_amp83 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=25e-6
m2 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=93e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=600e-6
m4 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
m5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=218e-6
m6 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=218e-6
m7 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=25e-6
m8 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=35e-6
m9 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=93e-6
m10 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos4 L=2e-6 W=19e-6
m11 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=35e-6
m12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=600e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=25e-6
m14 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=6e-6 W=129e-6
m15 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=6e-6 W=129e-6
m16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=197e-6
m17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=197e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp83

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 2.36101 mW
** Area: 11034 (mu_m)^2
** Transit frequency: 3.01801 MHz
** Transit frequency with error factor: 3.01768 MHz
** Slew rate: 10.6582 V/mu_s
** Phase margin: 79.6412°
** CMRR: 134 dB
** negPSRR: 37 dB
** posPSRR: 32 dB
** VoutMax: 4.30001 V
** VoutMin: 0.930001 V
** VcmMax: 4.67001 V
** VcmMin: 1.71001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00551e+07 muA
** DiodeTransistorPmos: -1.19233e+08 muA
** DiodeTransistorPmos: -1.19233e+08 muA
** NormalTransistorNmos: 2.38466e+08 muA
** DiodeTransistorNmos: 2.38465e+08 muA
** NormalTransistorNmos: 1.19234e+08 muA
** NormalTransistorNmos: 1.19234e+08 muA
** NormalTransistorNmos: 1.06744e+08 muA
** DiodeTransistorNmos: 1.06743e+08 muA
** NormalTransistorPmos: -1.06743e+08 muA
** NormalTransistorPmos: -1.06744e+08 muA
** NormalTransistorNmos: 1.06939e+08 muA
** NormalTransistorPmos: -1.06938e+08 muA
** NormalTransistorPmos: -1.06939e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.00559e+07 muA


** Expected Voltages: 
** ibias: 1.14501  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 4.26101  V
** inStageBiasComplementarySecondStage: 0.569001  V
** innerComplementarySecondStage: 1.33701  V
** out: 2.5  V
** outFirstStage: 4.26101  V
** outSourceVoltageBiasXXnXX1: 0.573001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.52501  V
** innerTransconductance: 4.77501  V
** inner: 4.77501  V
** inner: 0.571001  V


.END