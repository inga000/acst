** Name: two_stage_single_output_op_amp_55_9

.MACRO two_stage_single_output_op_amp_55_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=10e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=7e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=410e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=6e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=28e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=28e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=9e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=410e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=42e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=36e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=36e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=210e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=42e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=18e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_55_9

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 5.88401 mW
** Area: 6109 (mu_m)^2
** Transit frequency: 5.44601 MHz
** Transit frequency with error factor: 5.44555 MHz
** Slew rate: 4.73946 V/mu_s
** Phase margin: 64.1713°
** CMRR: 144 dB
** VoutMax: 4.25 V
** VoutMin: 1.25 V
** VcmMax: 5.17001 V
** VcmMin: 1.05001 V


** Expected Currents: 
** NormalTransistorPmos: -1.79349e+07 muA
** NormalTransistorPmos: -2.02769e+07 muA
** NormalTransistorPmos: -2.13969e+07 muA
** NormalTransistorPmos: -3.64989e+07 muA
** NormalTransistorPmos: -2.13969e+07 muA
** NormalTransistorPmos: -3.64989e+07 muA
** DiodeTransistorNmos: 2.13961e+07 muA
** NormalTransistorNmos: 2.13951e+07 muA
** NormalTransistorNmos: 2.13961e+07 muA
** DiodeTransistorNmos: 2.13951e+07 muA
** NormalTransistorNmos: 3.02011e+07 muA
** NormalTransistorNmos: 1.51011e+07 muA
** NormalTransistorNmos: 1.51011e+07 muA
** NormalTransistorNmos: 1.04566e+09 muA
** DiodeTransistorNmos: 1.04566e+09 muA
** NormalTransistorPmos: -1.04565e+09 muA
** DiodeTransistorNmos: 1.79341e+07 muA
** NormalTransistorNmos: 1.79331e+07 muA
** DiodeTransistorNmos: 2.02761e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.65801  V
** outSourceVoltageBiasXXnXX1: 0.829001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.850001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.629001  V
** innerTransistorStack1Load2: 0.629001  V
** out1: 1.19301  V
** sourceGCC1: 4.13001  V
** sourceGCC2: 4.13001  V
** sourceTransconductance: 1.89901  V
** inner: 0.825001  V


.END