.suckt  symmetrical_op_amp86 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_MainBias_1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_3 out2FirstStage out2FirstStage out1FirstStage out1FirstStage nmos
m_Symmetrical_FirstStage_Load_4 out1FirstStage out1FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Load_5 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage nmos
m_Symmetrical_FirstStage_Load_6 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_StageBias_7 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Transconductor_8 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_Symmetrical_FirstStage_Transconductor_9 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_Transconductor_10 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_Symmetrical_SecondStage1_Transconductor_11 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_StageBias_12 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m_Symmetrical_SecondStage1_StageBias_13 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_14 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_15 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_17 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_18 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Symmetrical_MainBias_19 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp86

