** Name: two_stage_single_output_op_amp_73_9

.MACRO two_stage_single_output_op_amp_73_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=67e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=5e-6 W=23e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=11e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=58e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=113e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=37e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=24e-6
mFoldedCascodeFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=20e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=10e-6 W=67e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=16e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=7e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=58e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=10e-6 W=74e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=61e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=76e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=76e-6
mMainBias19 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=309e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=8e-6 W=509e-6
mFoldedCascodeFirstStageLoad21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=61e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=286e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_73_9

** Expected Performance Values: 
** Gain: 118 dB
** Power consumption: 4.82401 mW
** Area: 11495 (mu_m)^2
** Transit frequency: 2.95301 MHz
** Transit frequency with error factor: 2.95286 MHz
** Slew rate: 4.3345 V/mu_s
** Phase margin: 60.1606°
** CMRR: 137 dB
** VoutMax: 4.25 V
** VoutMin: 1.84001 V
** VcmMax: 5.10001 V
** VcmMin: 1.77001 V


** Expected Currents: 
** NormalTransistorPmos: -1.18158e+08 muA
** NormalTransistorPmos: -1.27955e+08 muA
** NormalTransistorPmos: -2.05149e+07 muA
** NormalTransistorPmos: -3.19029e+07 muA
** NormalTransistorPmos: -2.05149e+07 muA
** NormalTransistorPmos: -3.19029e+07 muA
** NormalTransistorNmos: 2.05141e+07 muA
** NormalTransistorNmos: 2.05141e+07 muA
** DiodeTransistorNmos: 2.05141e+07 muA
** NormalTransistorNmos: 2.27731e+07 muA
** NormalTransistorNmos: 2.27721e+07 muA
** NormalTransistorNmos: 1.13871e+07 muA
** NormalTransistorNmos: 1.13871e+07 muA
** NormalTransistorNmos: 6.34818e+08 muA
** DiodeTransistorNmos: 6.34817e+08 muA
** NormalTransistorPmos: -6.34817e+08 muA
** DiodeTransistorNmos: 1.18159e+08 muA
** NormalTransistorNmos: 1.1816e+08 muA
** DiodeTransistorNmos: 1.27956e+08 muA
** DiodeTransistorNmos: 1.27955e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.64001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 2.24201  V
** outSourceVoltageBiasXXnXX1: 1.12101  V
** outSourceVoltageBiasXXnXX2: 0.664001  V
** outSourceVoltageBiasXXpXX1: 4.13101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.595001  V
** innerStageBias: 0.795001  V
** out1: 1.18101  V
** sourceGCC1: 4.15901  V
** sourceGCC2: 4.15901  V
** sourceTransconductance: 1.83501  V
** inner: 1.12201  V


.END