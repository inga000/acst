** Name: two_stage_single_output_op_amp_5_1

.MACRO two_stage_single_output_op_amp_5_1 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=7e-6
m2 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=40e-6
m3 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=51e-6
m4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
m5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
m6 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=237e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=51e-6
m8 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=70e-6
m9 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=5e-6 W=128e-6
m10 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=36e-6
m11 out ibias sourcePmos sourcePmos pmos4 L=5e-6 W=599e-6
m12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=70e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_5_1

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 1.06601 mW
** Area: 5728 (mu_m)^2
** Transit frequency: 3.47301 MHz
** Transit frequency with error factor: 3.47018 MHz
** Slew rate: 3.5144 V/mu_s
** Phase margin: 60.1606°
** CMRR: 106 dB
** negPSRR: 107 dB
** posPSRR: 156 dB
** VoutMax: 4.74001 V
** VoutMin: 0.150001 V
** VcmMax: 4.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -8.97899e+06 muA
** NormalTransistorNmos: 1.62241e+07 muA
** NormalTransistorNmos: 1.62231e+07 muA
** NormalTransistorNmos: 1.62241e+07 muA
** NormalTransistorNmos: 1.62231e+07 muA
** NormalTransistorPmos: -3.24499e+07 muA
** NormalTransistorPmos: -1.62249e+07 muA
** NormalTransistorPmos: -1.62249e+07 muA
** NormalTransistorNmos: 1.5175e+08 muA
** NormalTransistorPmos: -1.5175e+08 muA
** DiodeTransistorNmos: 8.97801e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.22501  V


.END