** Name: two_stage_single_output_op_amp_61_3

.MACRO two_stage_single_output_op_amp_61_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=8e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=181e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=61e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=12e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=60e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=60e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=46e-6
mFoldedCascodeFirstStageLoad10 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=12e-6
mMainBias11 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=63e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=107e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=181e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=76e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=76e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=69e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=541e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=541e-6
mFoldedCascodeFirstStageLoad20 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=53e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.80001e-12
.EOM two_stage_single_output_op_amp_61_3

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 2.99501 mW
** Area: 7853 (mu_m)^2
** Transit frequency: 3.36901 MHz
** Transit frequency with error factor: 3.36892 MHz
** Slew rate: 3.95022 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 4.48001 V
** VoutMin: 0.590001 V
** VcmMax: 3.29001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.99981e+07 muA
** NormalTransistorNmos: 5.13711e+07 muA
** NormalTransistorNmos: 1.90151e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** NormalTransistorNmos: 1.90151e+07 muA
** NormalTransistorNmos: 2.85701e+07 muA
** DiodeTransistorPmos: -1.90159e+07 muA
** NormalTransistorPmos: -1.90159e+07 muA
** NormalTransistorPmos: -1.90159e+07 muA
** NormalTransistorPmos: -1.91129e+07 muA
** NormalTransistorPmos: -1.91139e+07 muA
** NormalTransistorPmos: -9.55599e+06 muA
** NormalTransistorPmos: -9.55599e+06 muA
** NormalTransistorNmos: 4.50388e+08 muA
** NormalTransistorPmos: -4.50387e+08 muA
** NormalTransistorPmos: -4.50388e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -2.99989e+07 muA
** DiodeTransistorPmos: -5.13719e+07 muA


** Expected Voltages: 
** ibias: 1.20201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.997001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.22001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.42601  V
** innerTransistorStack2Load2: 4.45001  V
** out1: 4.19301  V
** sourceGCC1: 0.522001  V
** sourceGCC2: 0.522001  V
** sourceTransconductance: 3.25101  V
** innerStageBias: 4.55401  V


.END