** Name: two_stage_single_output_op_amp_47_1

.MACRO two_stage_single_output_op_amp_47_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=7e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=5e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=64e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=64e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=186e-6
mFoldedCascodeFirstStageLoad9 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=15e-6
mMainBias10 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=14e-6
mMainBias11 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=36e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=172e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=68e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=68e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=190e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=190e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=485e-6
mFoldedCascodeFirstStageLoad19 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=172e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_47_1

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 5.82401 mW
** Area: 7810 (mu_m)^2
** Transit frequency: 4.83201 MHz
** Transit frequency with error factor: 4.8324 MHz
** Slew rate: 6.15101 V/mu_s
** Phase margin: 71.0468°
** CMRR: 142 dB
** VoutMax: 4.65001 V
** VoutMin: 0.580001 V
** VcmMax: 3.89001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 9.25201e+06 muA
** NormalTransistorNmos: 2.39061e+07 muA
** NormalTransistorNmos: 2.78951e+07 muA
** NormalTransistorNmos: 4.18551e+07 muA
** NormalTransistorNmos: 2.78951e+07 muA
** NormalTransistorNmos: 4.18551e+07 muA
** NormalTransistorPmos: -2.78959e+07 muA
** NormalTransistorPmos: -2.78969e+07 muA
** NormalTransistorPmos: -2.78959e+07 muA
** NormalTransistorPmos: -2.78969e+07 muA
** NormalTransistorPmos: -2.79229e+07 muA
** NormalTransistorPmos: -1.39609e+07 muA
** NormalTransistorPmos: -1.39609e+07 muA
** NormalTransistorNmos: 1.03801e+09 muA
** NormalTransistorPmos: -1.038e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.25299e+06 muA
** DiodeTransistorPmos: -2.39069e+07 muA


** Expected Voltages: 
** ibias: 1.18701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.982001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.72001  V
** outVoltageBiasXXpXX2: 4.08901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.28401  V
** innerTransistorStack1Load2: 4.49601  V
** innerTransistorStack2Load2: 4.49601  V
** sourceGCC1: 0.524001  V
** sourceGCC2: 0.524001  V
** sourceTransconductance: 3.26601  V


.END