.suckt  complementary_op_amp18 ibias in1 in2 out sourceNmos sourcePmos
m_Complementary_MainBias_1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m_Complementary_FirstStage_Load_3 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_4 out FirstStageYout1 FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos pmos
m_Complementary_FirstStage_Load_5 FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m_Complementary_FirstStage_Load_7 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_8 out FirstStageYout1 FirstStageYinnerSourceLoadNmos FirstStageYinnerSourceLoadNmos nmos
m_Complementary_FirstStage_Load_9 FirstStageYinnerSourceLoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_10 FirstStageYsourceTransconductanceNmos outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_Complementary_FirstStage_StageBias_11 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_12 FirstStageYsourceTransconductancePmos ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_Complementary_FirstStage_StageBias_13 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Transconductor_14 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_15 FirstStageYinnerSourceLoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_16 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m_Complementary_FirstStage_Transconductor_17 FirstStageYinnerSourceLoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c_Complementary_Load_Capacitor_1 out sourceNmos 
m_Complementary_MainBias_18 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_Complementary_MainBias_19 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_MainBias_20 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_Complementary_MainBias_21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end complementary_op_amp18

