.suckt  two_stage_single_output_op_amp_34_8 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_3 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_5 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_SingleOutput_FirstStage_Load_6 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_StageBias_7 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_SingleOutput_FirstStage_StageBias_8 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Transconductor_9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_SingleOutput_FirstStage_Transconductor_10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_StageBias_11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m_SingleOutput_SecondStage1_StageBias_12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_Transconductor_13 out outFirstStage sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_14 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_SingleOutput_MainBias_15 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_16 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m_SingleOutput_MainBias_17 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_18 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_19 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_34_8

