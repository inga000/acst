.suckt  two_stage_fully_differential_op_amp_41_9 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m4 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m5 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m6 outFeedback outFeedback sourceNmos sourceNmos nmos
m7 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m8 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m9 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m11 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m13 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m14 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m15 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m16 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m17 sourceTransconductance outVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m18 FirstStageYinnerStageBias inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m19 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m20 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m21 out1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m22 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m23 out1 out1FirstStage sourcePmos sourcePmos pmos
m24 out2 ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m25 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m26 out2 out2FirstStage sourcePmos sourcePmos pmos
m27 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m28 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m29 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
m30 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m31 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
m32 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m33 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_41_9

