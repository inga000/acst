** Name: two_stage_single_output_op_amp_79_10

.MACRO two_stage_single_output_op_amp_79_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=10e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
mMainBias4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=63e-6
mFoldedCascodeFirstStageStageBias5 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=55e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=52e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=52e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=63e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=101e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=101e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=79e-6
mMainBias12 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=165e-6
mSecondStage1StageBias13 out ibias sourceNmos sourceNmos nmos4 L=9e-6 W=600e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=63e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=13e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=129e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=390e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=390e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=570e-6
mMainBias20 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=204e-6
mSecondStage1Transconductor21 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=579e-6
mFoldedCascodeFirstStageLoad22 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=129e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.30001e-12
.EOM two_stage_single_output_op_amp_79_10

** Expected Performance Values: 
** Gain: 139 dB
** Power consumption: 4.94001 mW
** Area: 14186 (mu_m)^2
** Transit frequency: 7.93001 MHz
** Transit frequency with error factor: 7.92982 MHz
** Slew rate: 7.12399 V/mu_s
** Phase margin: 60.1606°
** CMRR: 142 dB
** VoutMax: 4.52001 V
** VoutMin: 0.320001 V
** VcmMax: 5.25 V
** VcmMin: 1.47001 V


** Expected Currents: 
** NormalTransistorNmos: 1.62454e+08 muA
** NormalTransistorNmos: 1.30451e+07 muA
** NormalTransistorPmos: -4.17759e+07 muA
** NormalTransistorPmos: -5.23909e+07 muA
** NormalTransistorPmos: -7.98739e+07 muA
** NormalTransistorPmos: -5.23909e+07 muA
** NormalTransistorPmos: -7.98739e+07 muA
** NormalTransistorNmos: 5.23901e+07 muA
** NormalTransistorNmos: 5.23891e+07 muA
** NormalTransistorNmos: 5.23901e+07 muA
** NormalTransistorNmos: 5.23891e+07 muA
** NormalTransistorNmos: 5.49631e+07 muA
** NormalTransistorNmos: 5.49621e+07 muA
** NormalTransistorNmos: 2.74821e+07 muA
** NormalTransistorNmos: 2.74821e+07 muA
** NormalTransistorNmos: 6.01015e+08 muA
** NormalTransistorPmos: -6.01014e+08 muA
** NormalTransistorPmos: -6.01015e+08 muA
** DiodeTransistorNmos: 4.17751e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.62453e+08 muA
** DiodeTransistorPmos: -1.30459e+07 muA


** Expected Voltages: 
** ibias: 0.730001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11101  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.19201  V
** outVoltageBiasXXpXX2: 4.28401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.525001  V
** innerTransistorStack1Load2: 0.507001  V
** innerTransistorStack2Load2: 0.508001  V
** out1: 0.713001  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.49001  V


.END