.suckt  complementary_op_amp15 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m5 FirstStageYinnerTransistorStack1LoadPmos FirstStageYout1 sourcePmos sourcePmos pmos
m6 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m7 FirstStageYinnerTransistorStack2LoadPmos FirstStageYout1 sourcePmos sourcePmos pmos
m8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m9 FirstStageYinnerTransistorStack1LoadNmos FirstStageYout1 sourceNmos sourceNmos nmos
m10 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m11 FirstStageYinnerTransistorStack2LoadNmos FirstStageYout1 sourceNmos sourceNmos nmos
m12 FirstStageYsourceTransconductanceNmos outVoltageBiasXXnXX1 FirstStageYinnerStageBiasNmos FirstStageYinnerStageBiasNmos nmos
m13 FirstStageYinnerStageBiasNmos inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m14 FirstStageYsourceTransconductancePmos outVoltageBiasXXpXX1 FirstStageYinnerStageBiasPmos FirstStageYinnerStageBiasPmos pmos
m15 FirstStageYinnerStageBiasPmos ibias sourcePmos sourcePmos pmos
m16 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m17 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m18 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m19 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c1 out sourceNmos 
m20 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m21 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m22 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m23 ibias ibias sourcePmos sourcePmos pmos
.end complementary_op_amp15

