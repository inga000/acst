** Name: two_stage_single_output_op_amp_53_5

.MACRO two_stage_single_output_op_amp_53_5 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=14e-6
m2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=56e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=59e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=52e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=582e-6
m7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=63e-6
m8 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=423e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=260e-6
m10 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=56e-6
m11 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=136e-6
m12 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
m13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=24e-6
m14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=24e-6
m15 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=77e-6
m16 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=582e-6
m17 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=19e-6
m18 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=19e-6
m19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
m20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
m21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=52e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.70001e-12
.EOM two_stage_single_output_op_amp_53_5

** Expected Performance Values: 
** Gain: 117 dB
** Power consumption: 8.08001 mW
** Area: 11844 (mu_m)^2
** Transit frequency: 6.40001 MHz
** Transit frequency with error factor: 6.4003 MHz
** Slew rate: 7.92835 V/mu_s
** Phase margin: 60.1606°
** CMRR: 136 dB
** VoutMax: 3.01001 V
** VoutMin: 0.620001 V
** VcmMax: 4.68001 V
** VcmMin: 0.790001 V


** Expected Currents: 
** NormalTransistorNmos: 9.54311e+07 muA
** NormalTransistorNmos: 2.99525e+08 muA
** NormalTransistorPmos: -5.33309e+07 muA
** NormalTransistorPmos: -8.03469e+07 muA
** NormalTransistorPmos: -5.33309e+07 muA
** NormalTransistorPmos: -8.03469e+07 muA
** DiodeTransistorNmos: 5.33301e+07 muA
** DiodeTransistorNmos: 5.33291e+07 muA
** NormalTransistorNmos: 5.33301e+07 muA
** NormalTransistorNmos: 5.33291e+07 muA
** NormalTransistorNmos: 5.40311e+07 muA
** NormalTransistorNmos: 2.70151e+07 muA
** NormalTransistorNmos: 2.70151e+07 muA
** NormalTransistorNmos: 1.05045e+09 muA
** NormalTransistorPmos: -1.05044e+09 muA
** DiodeTransistorPmos: -1.05044e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.54319e+07 muA
** NormalTransistorPmos: -9.54329e+07 muA
** DiodeTransistorPmos: -2.99524e+08 muA
** DiodeTransistorPmos: -2.99525e+08 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 2.39201  V
** out: 2.5  V
** outFirstStage: 1.02601  V
** outInputVoltageBiasXXpXX1: 2.44401  V
** outSourceVoltageBiasXXpXX1: 3.72201  V
** outSourceVoltageBiasXXpXX2: 3.70601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.676001  V
** innerTransistorStack2Load2: 0.676001  V
** out1: 1.23101  V
** sourceGCC1: 3.51401  V
** sourceGCC2: 3.51401  V
** sourceTransconductance: 1.89501  V
** inner: 3.72101  V


.END