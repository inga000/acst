** Name: symmetrical_op_amp13

.MACRO symmetrical_op_amp13 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=26e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=26e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=20e-6
mSecondStage1StageBias5 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=29e-6
mSecondStage1Transconductor6 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=48e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor7 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=48e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=4e-6 W=22e-6
mSecondStage1Transconductor9 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=22e-6
mSymmetricalFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=80e-6
mMainBias11 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=3e-6 W=37e-6
mSymmetricalFirstStageTransconductor12 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=150e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias13 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=29e-6
mSecondStage1StageBias14 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=1e-6 W=85e-6
mSymmetricalFirstStageTransconductor15 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=150e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp13

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 0.769001 mW
** Area: 2770 (mu_m)^2
** Transit frequency: 3.42901 MHz
** Transit frequency with error factor: 3.42945 MHz
** Slew rate: 3.70296 V/mu_s
** Phase margin: 80.7871°
** CMRR: 149 dB
** negPSRR: 50 dB
** posPSRR: 59 dB
** VoutMax: 3.68001 V
** VoutMin: 0.470001 V
** VcmMax: 3.97001 V
** VcmMin: 0.0300001 V


** Expected Currents: 
** NormalTransistorPmos: -1.88509e+07 muA
** DiodeTransistorNmos: 2.03791e+07 muA
** DiodeTransistorNmos: 2.03791e+07 muA
** NormalTransistorPmos: -4.07599e+07 muA
** NormalTransistorPmos: -2.03799e+07 muA
** NormalTransistorPmos: -2.03799e+07 muA
** NormalTransistorNmos: 3.70751e+07 muA
** NormalTransistorNmos: 3.70761e+07 muA
** NormalTransistorPmos: -3.70759e+07 muA
** DiodeTransistorPmos: -3.70769e+07 muA
** NormalTransistorPmos: -3.70779e+07 muA
** NormalTransistorNmos: 3.70771e+07 muA
** NormalTransistorNmos: 3.70761e+07 muA
** DiodeTransistorNmos: 1.88501e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.14501  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.878001  V
** inSourceTransconductanceComplementarySecondStage: 0.597001  V
** inStageBiasComplementarySecondStage: 3.83501  V
** innerComplementarySecondStage: 3.11401  V
** out: 2.5  V
** outFirstStage: 0.597001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.23801  V
** innerTransconductance: 0.192001  V
** inner: 0.192001  V


.END