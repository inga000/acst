.suckt  two_stage_fully_differential_op_amp_16_12 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_3 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_4 outInputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_5 outVoltageBiasXXnXX3 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_6 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_7 outFeedback outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_8 FeedbackStageYsourceTransconductance1 outVoltageBiasXXnXX3 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYinnerStageBias1 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_10 FeedbackStageYsourceTransconductance2 outVoltageBiasXXnXX3 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m_FullyDifferential_FeedbackdStage_StageBias_11 FeedbackStageYinnerStageBias2 ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackStage_Transconductor_12 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_13 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_14 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FeedbackStage_Transconductor_15 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FirstStage_Load_16 out1FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m_FullyDifferential_FirstStage_Load_17 FirstStageYinnerTransistorStack1Load1 outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_18 out2FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_FullyDifferential_FirstStage_Load_19 FirstStageYinnerTransistorStack2Load1 outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_StageBias_20 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Transconductor_21 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_FullyDifferential_FirstStage_Transconductor_22 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_StageBias_23 out1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_FullyDifferential_SecondStage1_StageBias_24 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_Transconductor_25 out1 outVoltageBiasXXpXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
m_FullyDifferential_SecondStage1_Transconductor_26 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_StageBias_27 out2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m_FullyDifferential_SecondStage2_StageBias_28 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_Transconductor_29 out2 outVoltageBiasXXpXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
m_FullyDifferential_SecondStage2_Transconductor_30 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_31 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_FullyDifferential_MainBias_32 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_33 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
m_FullyDifferential_MainBias_34 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_35 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_36 ibias ibias sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_37 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_38 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_16_12

