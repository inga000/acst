** Name: two_stage_single_output_op_amp_60_9

.MACRO two_stage_single_output_op_amp_60_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=74e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=15e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=562e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=61e-6
m5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=85e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=216e-6
m7 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=52e-6
m8 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=562e-6
m9 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=40e-6
m10 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=40e-6
m11 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=54e-6
m12 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=54e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=15e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=494e-6
m15 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=301e-6
m16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=5e-6 W=114e-6
m17 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=284e-6
m18 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=52e-6
m19 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=16e-6
m20 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=16e-6
m21 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=216e-6
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=85e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_60_9

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 6.91301 mW
** Area: 12562 (mu_m)^2
** Transit frequency: 4.25101 MHz
** Transit frequency with error factor: 4.25064 MHz
** Slew rate: 4.19346 V/mu_s
** Phase margin: 69.328°
** CMRR: 141 dB
** VoutMax: 4.25 V
** VoutMin: 0.730001 V
** VcmMax: 3.26001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorPmos: -3.32469e+07 muA
** NormalTransistorPmos: -3.56459e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 3.19131e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 3.19131e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** DiodeTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -2.57339e+07 muA
** DiodeTransistorPmos: -2.57329e+07 muA
** NormalTransistorPmos: -1.28669e+07 muA
** NormalTransistorPmos: -1.28669e+07 muA
** NormalTransistorNmos: 1.22988e+09 muA
** DiodeTransistorNmos: 1.22988e+09 muA
** NormalTransistorPmos: -1.22987e+09 muA
** DiodeTransistorNmos: 3.32461e+07 muA
** NormalTransistorNmos: 3.32451e+07 muA
** DiodeTransistorNmos: 3.56451e+07 muA
** DiodeTransistorNmos: 3.56461e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.12801  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.13101  V
** outSourceVoltageBiasXXnXX1: 0.566001  V
** outSourceVoltageBiasXXnXX2: 0.572001  V
** outSourceVoltageBiasXXpXX1: 4.23701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.14901  V
** out1: 3.36801  V
** sourceGCC1: 0.573001  V
** sourceGCC2: 0.573001  V
** sourceTransconductance: 3.27601  V
** inner: 0.564001  V
** inner: 4.23401  V


.END