** Name: two_stage_single_output_op_amp_51_9

.MACRO two_stage_single_output_op_amp_51_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=47e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=13e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=223e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=34e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=24e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=47e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=13e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=13e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=13e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=223e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=13e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=128e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=54e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=54e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=539e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=128e-6
mMainBias19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=110e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=48e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_51_9

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 5.30501 mW
** Area: 9893 (mu_m)^2
** Transit frequency: 3.46301 MHz
** Transit frequency with error factor: 3.46274 MHz
** Slew rate: 3.81467 V/mu_s
** Phase margin: 62.4525°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 1.64001 V
** VcmMax: 5.12001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorPmos: -5.32399e+07 muA
** NormalTransistorPmos: -2.32579e+07 muA
** NormalTransistorPmos: -1.73279e+07 muA
** NormalTransistorPmos: -2.62049e+07 muA
** NormalTransistorPmos: -1.73279e+07 muA
** NormalTransistorPmos: -2.62049e+07 muA
** NormalTransistorNmos: 1.73271e+07 muA
** NormalTransistorNmos: 1.73271e+07 muA
** DiodeTransistorNmos: 1.73271e+07 muA
** NormalTransistorNmos: 1.77511e+07 muA
** NormalTransistorNmos: 8.87601e+06 muA
** NormalTransistorNmos: 8.87601e+06 muA
** NormalTransistorNmos: 9.12114e+08 muA
** DiodeTransistorNmos: 9.12113e+08 muA
** NormalTransistorPmos: -9.12113e+08 muA
** DiodeTransistorNmos: 5.32391e+07 muA
** NormalTransistorNmos: 5.32381e+07 muA
** DiodeTransistorNmos: 2.32571e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 2.04801  V
** outSourceVoltageBiasXXnXX1: 1.02401  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** outVoltageBiasXXnXX2: 0.605001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.591001  V
** out1: 1.17301  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.91501  V
** inner: 1.01801  V


.END