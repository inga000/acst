** Name: two_stage_single_output_op_amp_15_2

.MACRO two_stage_single_output_op_amp_15_2 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=33e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mSecondStage1StageBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=28e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=49e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=46e-6
mSecondStage1Transconductor6 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=327e-6
mMainBias7 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=479e-6
mSecondStage1Transconductor8 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=110e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=33e-6
mSimpleFirstStageStageBias10 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=78e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=3e-6 W=51e-6
mSecondStage1StageBias13 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=478e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=10e-6
mMainBias15 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=48e-6
mMainBias16 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=460e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_15_2

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 1.84001 mW
** Area: 9832 (mu_m)^2
** Transit frequency: 2.64901 MHz
** Transit frequency with error factor: 2.64422 MHz
** Slew rate: 3.50007 V/mu_s
** Phase margin: 60.7336°
** CMRR: 97 dB
** negPSRR: 98 dB
** posPSRR: 122 dB
** VoutMax: 4.85001 V
** VoutMin: 0.350001 V
** VcmMax: 3.28001 V
** VcmMin: 0.0100001 V


** Expected Currents: 
** NormalTransistorNmos: 1.30332e+08 muA
** NormalTransistorPmos: -9.87599e+06 muA
** NormalTransistorPmos: -9.36489e+07 muA
** DiodeTransistorNmos: 7.89801e+06 muA
** NormalTransistorNmos: 7.89801e+06 muA
** NormalTransistorPmos: -1.57989e+07 muA
** NormalTransistorPmos: -1.57999e+07 muA
** NormalTransistorPmos: -7.89899e+06 muA
** NormalTransistorPmos: -7.89899e+06 muA
** NormalTransistorNmos: 9.83641e+07 muA
** NormalTransistorNmos: 9.83631e+07 muA
** NormalTransistorPmos: -9.83649e+07 muA
** DiodeTransistorNmos: 9.87501e+06 muA
** DiodeTransistorNmos: 9.36481e+07 muA
** DiodeTransistorPmos: -1.30331e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.74301  V
** out: 2.5  V
** outFirstStage: 0.573001  V
** outVoltageBiasXXnXX0: 0.555001  V
** outVoltageBiasXXnXX1: 0.751001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.53401  V
** out1: 0.573001  V
** sourceTransconductance: 3.27401  V
** innerTransconductance: 0.168001  V


.END