** Name: two_stage_single_output_op_amp_48_8

.MACRO two_stage_single_output_op_amp_48_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=23e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=140e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=140e-6
mMainBias5 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=89e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 outInputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=18e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=37e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=37e-6
mSecondStage1StageBias9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=521e-6
mSecondStage1StageBias10 out outInputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=446e-6
mFoldedCascodeFirstStageLoad11 outFirstStage outInputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=18e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=6e-6 W=140e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=198e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=198e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=414e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=98e-6
mFoldedCascodeFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=2e-6 W=140e-6
mMainBias18 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=407e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_48_8

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 6.00801 mW
** Area: 10902 (mu_m)^2
** Transit frequency: 4.50501 MHz
** Transit frequency with error factor: 4.50512 MHz
** Slew rate: 5.11591 V/mu_s
** Phase margin: 60.1606°
** CMRR: 143 dB
** VoutMax: 4.25 V
** VoutMin: 0.720001 V
** VcmMax: 4.06001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -4.57119e+07 muA
** NormalTransistorNmos: 4.67911e+07 muA
** NormalTransistorNmos: 7.04721e+07 muA
** NormalTransistorNmos: 4.67911e+07 muA
** NormalTransistorNmos: 7.04721e+07 muA
** DiodeTransistorPmos: -4.67919e+07 muA
** NormalTransistorPmos: -4.67929e+07 muA
** NormalTransistorPmos: -4.67919e+07 muA
** DiodeTransistorPmos: -4.67929e+07 muA
** NormalTransistorPmos: -4.73589e+07 muA
** NormalTransistorPmos: -2.36799e+07 muA
** NormalTransistorPmos: -2.36799e+07 muA
** NormalTransistorNmos: 9.95034e+08 muA
** NormalTransistorNmos: 9.95033e+08 muA
** NormalTransistorPmos: -9.95033e+08 muA
** DiodeTransistorNmos: 4.57111e+07 muA
** DiodeTransistorNmos: 4.57121e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.11301  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.10001  V
** innerTransistorStack1Load2: 4.09901  V
** out1: 3.34201  V
** sourceGCC1: 0.532001  V
** sourceGCC2: 0.532001  V
** sourceTransconductance: 3.24701  V
** innerStageBias: 0.545001  V


.END