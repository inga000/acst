** Name: two_stage_single_output_op_amp_52_10

.MACRO two_stage_single_output_op_amp_52_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=188e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=49e-6
m5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=506e-6
m6 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=177e-6
m7 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=423e-6
m8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=6e-6
m9 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=77e-6
m10 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=10e-6 W=188e-6
m11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=50e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=50e-6
m13 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=26e-6
m14 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=539e-6
m15 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=414e-6
m16 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=70e-6
m17 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=70e-6
m18 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=257e-6
m19 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=257e-6
m20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=562e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 7.10001e-12
.EOM two_stage_single_output_op_amp_52_10

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 5.97901 mW
** Area: 13519 (mu_m)^2
** Transit frequency: 5.06701 MHz
** Transit frequency with error factor: 5.06694 MHz
** Slew rate: 5.11717 V/mu_s
** Phase margin: 60.1606°
** CMRR: 144 dB
** VoutMax: 4.25 V
** VoutMin: 0.220001 V
** VcmMax: 5.22001 V
** VcmMin: 0.790001 V


** Expected Currents: 
** NormalTransistorNmos: 2.48758e+08 muA
** NormalTransistorNmos: 1.07939e+08 muA
** NormalTransistorPmos: -1.15844e+08 muA
** NormalTransistorPmos: -3.64469e+07 muA
** NormalTransistorPmos: -5.46689e+07 muA
** NormalTransistorPmos: -3.64499e+07 muA
** NormalTransistorPmos: -5.46739e+07 muA
** DiodeTransistorNmos: 3.64481e+07 muA
** NormalTransistorNmos: 3.64491e+07 muA
** NormalTransistorNmos: 3.64481e+07 muA
** NormalTransistorNmos: 3.64471e+07 muA
** NormalTransistorNmos: 1.82231e+07 muA
** NormalTransistorNmos: 1.82231e+07 muA
** NormalTransistorNmos: 6.03825e+08 muA
** NormalTransistorPmos: -6.03824e+08 muA
** NormalTransistorPmos: -6.03825e+08 muA
** DiodeTransistorNmos: 1.15845e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.48757e+08 muA
** DiodeTransistorPmos: -1.07938e+08 muA


** Expected Voltages: 
** ibias: 0.629001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.14201  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.08801  V
** outVoltageBiasXXpXX2: 4.24701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.357001  V
** out1: 0.556001  V
** sourceGCC1: 4.49101  V
** sourceGCC2: 4.49101  V
** sourceTransconductance: 1.93401  V
** innerTransconductance: 4.65201  V


.END