** Name: two_stage_single_output_op_amp_152_9

.MACRO two_stage_single_output_op_amp_152_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=6e-6 W=34e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=34e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=36e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=509e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=143e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageTransconductor8 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=39e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=10e-6 W=34e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=154e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=36e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=509e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=6e-6 W=34e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=39e-6
mSimpleFirstStageLoad15 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=264e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=166e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=166e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=376e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=264e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=88e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.80001e-12
.EOM two_stage_single_output_op_amp_152_9

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 8.71901 mW
** Area: 7368 (mu_m)^2
** Transit frequency: 5.60001 MHz
** Transit frequency with error factor: 5.59687 MHz
** Slew rate: 5.52774 V/mu_s
** Phase margin: 60.1606°
** CMRR: 116 dB
** VoutMax: 4.25 V
** VoutMin: 0.75 V
** VcmMax: 4.98001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorPmos: -8.92209e+07 muA
** NormalTransistorPmos: -3.04159e+07 muA
** DiodeTransistorNmos: 1.49471e+08 muA
** NormalTransistorNmos: 1.49472e+08 muA
** NormalTransistorNmos: 1.49473e+08 muA
** DiodeTransistorNmos: 1.49472e+08 muA
** NormalTransistorPmos: -1.65765e+08 muA
** NormalTransistorPmos: -1.65766e+08 muA
** NormalTransistorPmos: -1.65767e+08 muA
** NormalTransistorPmos: -1.65766e+08 muA
** NormalTransistorNmos: 3.25911e+07 muA
** NormalTransistorNmos: 1.62951e+07 muA
** NormalTransistorNmos: 1.62951e+07 muA
** NormalTransistorNmos: 1.27256e+09 muA
** DiodeTransistorNmos: 1.27256e+09 muA
** NormalTransistorPmos: -1.27255e+09 muA
** DiodeTransistorNmos: 8.92201e+07 muA
** NormalTransistorNmos: 8.92191e+07 muA
** DiodeTransistorNmos: 3.04151e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.15201  V
** outSourceVoltageBiasXXnXX1: 0.576001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerTransistorStack1Load1: 1.13001  V
** innerTransistorStack1Load2: 4.16001  V
** innerTransistorStack2Load1: 1.12901  V
** innerTransistorStack2Load2: 4.16001  V
** sourceTransconductance: 1.93801  V
** inner: 0.576001  V


.END