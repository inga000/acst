** Name: two_stage_single_output_op_amp_9_10

.MACRO two_stage_single_output_op_amp_9_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
m2 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
m3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=530e-6
m4 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=145e-6
m5 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=551e-6
m6 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=269e-6
m7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=145e-6
m8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=85e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=495e-6
m10 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
m11 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=5e-6 W=530e-6
m12 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=320e-6
Capacitor1 outFirstStage out 19.8001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_9_10

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 8.92901 mW
** Area: 14087 (mu_m)^2
** Transit frequency: 5.36801 MHz
** Transit frequency with error factor: 5.36379 MHz
** Slew rate: 8.33989 V/mu_s
** Phase margin: 60.1606°
** CMRR: 102 dB
** negPSRR: 109 dB
** posPSRR: 97 dB
** VoutMax: 4.25 V
** VoutMin: 0.260001 V
** VcmMax: 4.41001 V
** VcmMin: 0.920001 V


** Expected Currents: 
** NormalTransistorNmos: 5.27977e+08 muA
** NormalTransistorPmos: -8.33819e+07 muA
** NormalTransistorPmos: -8.33819e+07 muA
** DiodeTransistorPmos: -8.33819e+07 muA
** NormalTransistorNmos: 1.66763e+08 muA
** NormalTransistorNmos: 8.33811e+07 muA
** NormalTransistorNmos: 8.33811e+07 muA
** NormalTransistorNmos: 1.08101e+09 muA
** NormalTransistorPmos: -1.081e+09 muA
** NormalTransistorPmos: -1.081e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.27976e+08 muA


** Expected Voltages: 
** ibias: 0.670001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.00201  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.22601  V
** out1: 3.44401  V
** sourceTransconductance: 1.84701  V
** innerTransconductance: 4.56601  V


.END