** Name: two_stage_single_output_op_amp_75_8

.MACRO two_stage_single_output_op_amp_75_8 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=230e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=86e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m6 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=274e-6
m7 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=23e-6
m8 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
m9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=86e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=58e-6
m11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=58e-6
m12 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=20e-6
m13 SecondStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=512e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=516e-6
m15 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=62e-6
m16 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=327e-6
m17 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=579e-6
m18 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=62e-6
m19 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=76e-6
m20 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=76e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.70001e-12
.EOM two_stage_single_output_op_amp_75_8

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 11.9621 mW
** Area: 6664 (mu_m)^2
** Transit frequency: 6.61801 MHz
** Transit frequency with error factor: 6.61829 MHz
** Slew rate: 6.7253 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 4.25 V
** VoutMin: 0.410001 V
** VcmMax: 5.17001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorPmos: -3.31537e+08 muA
** NormalTransistorPmos: -5.76934e+08 muA
** NormalTransistorPmos: -4.52139e+07 muA
** NormalTransistorPmos: -7.70539e+07 muA
** NormalTransistorPmos: -4.52139e+07 muA
** NormalTransistorPmos: -7.70539e+07 muA
** DiodeTransistorNmos: 4.52131e+07 muA
** NormalTransistorNmos: 4.52131e+07 muA
** NormalTransistorNmos: 4.52131e+07 muA
** NormalTransistorNmos: 6.36771e+07 muA
** NormalTransistorNmos: 6.36761e+07 muA
** NormalTransistorNmos: 3.18391e+07 muA
** NormalTransistorNmos: 3.18391e+07 muA
** NormalTransistorNmos: 1.30979e+09 muA
** NormalTransistorNmos: 1.30979e+09 muA
** NormalTransistorPmos: -1.30978e+09 muA
** DiodeTransistorNmos: 3.31538e+08 muA
** DiodeTransistorNmos: 5.76935e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.02801  V
** outVoltageBiasXXnXX2: 0.578001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.429001  V
** innerTransistorStack2Load2: 0.470001  V
** out1: 0.627001  V
** sourceGCC1: 4.16301  V
** sourceGCC2: 4.16301  V
** sourceTransconductance: 1.86701  V
** innerStageBias: 0.385001  V


.END