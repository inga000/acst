** Name: two_stage_single_output_op_amp_46_2

.MACRO two_stage_single_output_op_amp_46_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=152e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
m4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=170e-6
m5 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=176e-6
m6 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=288e-6
m7 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=27e-6
m8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=27e-6
m9 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=520e-6
m10 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=520e-6
m11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=30e-6
m12 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=75e-6
m13 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=379e-6
m14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=176e-6
m15 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=238e-6
m16 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=170e-6
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=13e-6
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=13e-6
m19 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=178e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.70001e-12
.EOM two_stage_single_output_op_amp_46_2

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 3.01201 mW
** Area: 14062 (mu_m)^2
** Transit frequency: 2.73101 MHz
** Transit frequency with error factor: 2.73072 MHz
** Slew rate: 6.81185 V/mu_s
** Phase margin: 60.1606°
** CMRR: 128 dB
** VoutMax: 4.72001 V
** VoutMin: 0.420001 V
** VcmMax: 3.41001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.15498e+08 muA
** NormalTransistorPmos: -3.63969e+07 muA
** NormalTransistorNmos: 8.06111e+07 muA
** NormalTransistorNmos: 1.23802e+08 muA
** NormalTransistorNmos: 8.06091e+07 muA
** NormalTransistorNmos: 1.23802e+08 muA
** DiodeTransistorPmos: -8.06119e+07 muA
** DiodeTransistorPmos: -8.06109e+07 muA
** NormalTransistorPmos: -8.06099e+07 muA
** NormalTransistorPmos: -8.06109e+07 muA
** NormalTransistorPmos: -8.63819e+07 muA
** NormalTransistorPmos: -4.31909e+07 muA
** NormalTransistorPmos: -4.31909e+07 muA
** NormalTransistorNmos: 1.82846e+08 muA
** NormalTransistorNmos: 1.82845e+08 muA
** NormalTransistorPmos: -1.82845e+08 muA
** DiodeTransistorNmos: 1.15499e+08 muA
** DiodeTransistorNmos: 3.63961e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.15201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.674001  V
** outVoltageBiasXXnXX1: 1.07901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.27301  V
** innerTransistorStack2Load2: 4.27301  V
** out1: 3.54901  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.80801  V
** innerTransconductance: 0.524001  V


.END