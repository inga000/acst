** Name: two_stage_single_output_op_amp_58_2

.MACRO two_stage_single_output_op_amp_58_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=22e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=6e-6
m3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=164e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=277e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=496e-6
m7 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=215e-6
m8 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=294e-6
m9 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=294e-6
m10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=240e-6
m11 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=353e-6
m12 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=215e-6
m13 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=138e-6
m14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=76e-6
m15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=76e-6
m16 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=496e-6
m17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=277e-6
m18 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
m19 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=522e-6
m20 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=9e-6 W=164e-6
m21 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=58e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 12.3001e-12
.EOM two_stage_single_output_op_amp_58_2

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 3.15901 mW
** Area: 15000 (mu_m)^2
** Transit frequency: 2.94901 MHz
** Transit frequency with error factor: 2.94268 MHz
** Slew rate: 6.59315 V/mu_s
** Phase margin: 60.1606°
** CMRR: 85 dB
** VoutMax: 4.84001 V
** VoutMin: 0.350001 V
** VcmMax: 3.04001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 6.57101e+07 muA
** NormalTransistorPmos: -2.54779e+07 muA
** NormalTransistorPmos: -1.04769e+07 muA
** NormalTransistorNmos: 8.19011e+07 muA
** NormalTransistorNmos: 1.40404e+08 muA
** NormalTransistorNmos: 8.18991e+07 muA
** NormalTransistorNmos: 1.404e+08 muA
** DiodeTransistorPmos: -8.18999e+07 muA
** NormalTransistorPmos: -8.18999e+07 muA
** NormalTransistorPmos: -1.17002e+08 muA
** DiodeTransistorPmos: -1.17003e+08 muA
** NormalTransistorPmos: -5.85009e+07 muA
** NormalTransistorPmos: -5.85009e+07 muA
** NormalTransistorNmos: 2.29302e+08 muA
** NormalTransistorNmos: 2.29301e+08 muA
** NormalTransistorPmos: -2.29301e+08 muA
** DiodeTransistorNmos: 2.54771e+07 muA
** DiodeTransistorNmos: 1.04761e+07 muA
** DiodeTransistorPmos: -6.57109e+07 muA
** NormalTransistorPmos: -6.57119e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.28001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.54601  V
** outSourceVoltageBiasXXpXX1: 4.27301  V
** outVoltageBiasXXnXX1: 0.905001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.93201  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.57001  V
** innerTransconductance: 0.304001  V
** inner: 4.27301  V


.END