** Name: two_stage_single_output_op_amp_58_10

.MACRO two_stage_single_output_op_amp_58_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=35e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=179e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=23e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=294e-6
mSecondStage1StageBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=45e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=102e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=86e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=86e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=596e-6
mFoldedCascodeFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=102e-6
mMainBias12 outVoltageBiasXXpXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=219e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=116e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=116e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=294e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=420e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=23e-6
mSecondStage1Transconductor18 out outVoltageBiasXXpXX2 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad19 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=179e-6
mMainBias20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=155e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=165e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 18.2001e-12
.EOM two_stage_single_output_op_amp_58_10

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 11.1391 mW
** Area: 7391 (mu_m)^2
** Transit frequency: 6.39501 MHz
** Transit frequency with error factor: 6.38774 MHz
** Slew rate: 6.17072 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.25 V
** VoutMin: 0.160001 V
** VcmMax: 3.15001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.56903e+08 muA
** NormalTransistorPmos: -6.74679e+07 muA
** NormalTransistorPmos: -7.23069e+07 muA
** NormalTransistorNmos: 1.12709e+08 muA
** NormalTransistorNmos: 1.77667e+08 muA
** NormalTransistorNmos: 1.12709e+08 muA
** NormalTransistorNmos: 1.77667e+08 muA
** DiodeTransistorPmos: -1.12708e+08 muA
** NormalTransistorPmos: -1.12708e+08 muA
** NormalTransistorPmos: -1.29913e+08 muA
** DiodeTransistorPmos: -1.29912e+08 muA
** NormalTransistorPmos: -6.49569e+07 muA
** NormalTransistorPmos: -6.49569e+07 muA
** NormalTransistorNmos: 1.25584e+09 muA
** NormalTransistorPmos: -1.25583e+09 muA
** NormalTransistorPmos: -1.25583e+09 muA
** DiodeTransistorNmos: 6.74671e+07 muA
** DiodeTransistorNmos: 7.23061e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -4.56902e+08 muA


** Expected Voltages: 
** ibias: 3.32801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.02701  V
** outSourceVoltageBiasXXpXX1: 4.16501  V
** outVoltageBiasXXnXX1: 0.923001  V
** outVoltageBiasXXnXX2: 0.562001  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.01501  V
** sourceGCC1: 0.357001  V
** sourceGCC2: 0.357001  V
** sourceTransconductance: 3.24101  V
** innerTransconductance: 4.59101  V
** inner: 4.16101  V


.END