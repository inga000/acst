** Name: two_stage_single_output_op_amp_206_7

.MACRO two_stage_single_output_op_amp_206_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=17e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=17e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=143e-6
mSimpleFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=16e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=10e-6 W=17e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=31e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=15e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=143e-6
mSecondStage1StageBias12 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=488e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=7e-6 W=17e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=31e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=77e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=77e-6
mSimpleFirstStageLoad17 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=39e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=272e-6
mSimpleFirstStageLoad19 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=39e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=151e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=45e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_206_7

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 8.76801 mW
** Area: 7490 (mu_m)^2
** Transit frequency: 3.58601 MHz
** Transit frequency with error factor: 3.58508 MHz
** Slew rate: 3.5002 V/mu_s
** Phase margin: 72.1927°
** CMRR: 116 dB
** VoutMax: 4.25 V
** VoutMin: 0.480001 V
** VcmMax: 4.84001 V
** VcmMin: 1.51001 V


** Expected Currents: 
** NormalTransistorPmos: -1.51881e+08 muA
** NormalTransistorPmos: -4.54059e+07 muA
** DiodeTransistorNmos: 6.98151e+07 muA
** NormalTransistorNmos: 6.98161e+07 muA
** NormalTransistorNmos: 6.98151e+07 muA
** DiodeTransistorNmos: 6.98161e+07 muA
** NormalTransistorPmos: -7.77309e+07 muA
** NormalTransistorPmos: -7.77319e+07 muA
** NormalTransistorPmos: -7.77309e+07 muA
** NormalTransistorPmos: -7.77319e+07 muA
** NormalTransistorNmos: 1.58301e+07 muA
** DiodeTransistorNmos: 1.58291e+07 muA
** NormalTransistorNmos: 7.91501e+06 muA
** NormalTransistorNmos: 7.91501e+06 muA
** NormalTransistorNmos: 1.38087e+09 muA
** NormalTransistorPmos: -1.38086e+09 muA
** DiodeTransistorNmos: 1.51882e+08 muA
** NormalTransistorNmos: 1.51881e+08 muA
** DiodeTransistorNmos: 4.54051e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.35601  V
** outSourceVoltageBiasXXnXX1: 0.678001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.887001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.10501  V
** innerTransistorStack1Load1: 1.10501  V
** innerTransistorStack1Load2: 4.29501  V
** innerTransistorStack2Load2: 4.29501  V
** out1: 2.09501  V
** sourceTransconductance: 1.93901  V
** inner: 0.676001  V


.END