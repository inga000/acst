** Name: two_stage_single_output_op_amp_16_2

.MACRO two_stage_single_output_op_amp_16_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=16e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=31e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=18e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=103e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=206e-6
m7 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=398e-6
m8 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=31e-6
m9 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=35e-6
m10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=108e-6
m11 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=14e-6
m12 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=367e-6
m13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=88e-6
m14 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
m15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=88e-6
m16 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=206e-6
m17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=103e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_16_2

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 1.32101 mW
** Area: 8134 (mu_m)^2
** Transit frequency: 3.30601 MHz
** Transit frequency with error factor: 3.30263 MHz
** Slew rate: 3.72641 V/mu_s
** Phase margin: 71.6198°
** CMRR: 100 dB
** negPSRR: 101 dB
** posPSRR: 127 dB
** VoutMax: 4.75 V
** VoutMin: 0.310001 V
** VcmMax: 3.36001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 8.47201e+06 muA
** NormalTransistorPmos: -3.94799e+06 muA
** NormalTransistorPmos: -7.89699e+06 muA
** DiodeTransistorNmos: 8.43501e+06 muA
** NormalTransistorNmos: 8.43501e+06 muA
** NormalTransistorPmos: -1.68729e+07 muA
** DiodeTransistorPmos: -1.68739e+07 muA
** NormalTransistorPmos: -8.43599e+06 muA
** NormalTransistorPmos: -8.43599e+06 muA
** NormalTransistorNmos: 2.07016e+08 muA
** NormalTransistorNmos: 2.07015e+08 muA
** NormalTransistorPmos: -2.07015e+08 muA
** DiodeTransistorNmos: 3.94701e+06 muA
** DiodeTransistorNmos: 7.89601e+06 muA
** DiodeTransistorPmos: -8.47299e+06 muA
** NormalTransistorPmos: -8.47399e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.711001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.54001  V
** outSourceVoltageBiasXXpXX1: 4.27001  V
** outVoltageBiasXXnXX0: 0.557001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceTransconductance: 3.24301  V
** innerTransconductance: 0.150001  V
** inner: 4.27001  V


.END