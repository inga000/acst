** Name: one_stage_single_output_op_amp93

.MACRO one_stage_single_output_op_amp93 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=4e-6
m3 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
m4 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
m5 out outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=67e-6
m6 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
m7 sourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=58e-6
m8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=67e-6
m9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=67e-6
m10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=67e-6
m11 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=160e-6
m12 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m13 FirstStageYout1 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp93

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 0.625001 mW
** Area: 1591 (mu_m)^2
** Transit frequency: 4.49901 MHz
** Transit frequency with error factor: 4.49877 MHz
** Slew rate: 4.74907 V/mu_s
** Phase margin: 87.0896°
** CMRR: 151 dB
** VoutMax: 3.61001 V
** VoutMin: 0.5 V
** VcmMax: 3.86001 V
** VcmMin: 0.75 V


** Expected Currents: 
** NormalTransistorNmos: 1.97531e+07 muA
** NormalTransistorPmos: -1.02139e+07 muA
** NormalTransistorNmos: 4.25381e+07 muA
** NormalTransistorNmos: 4.25371e+07 muA
** NormalTransistorPmos: -4.25389e+07 muA
** NormalTransistorPmos: -4.25379e+07 muA
** DiodeTransistorPmos: -4.25389e+07 muA
** NormalTransistorNmos: 9.52881e+07 muA
** NormalTransistorNmos: 4.25371e+07 muA
** NormalTransistorNmos: 4.25371e+07 muA
** DiodeTransistorNmos: 1.02131e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.97539e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 4.19601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack2Load2: 3.82001  V
** out1: 3.04401  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END