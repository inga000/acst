** Name: two_stage_single_output_op_amp_195_8

.MACRO two_stage_single_output_op_amp_195_8 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=4e-6 W=12e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=19e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=76e-6
mSimpleFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=99e-6
mSimpleFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=13e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=25e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=94e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mMainBias11 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=80e-6
mSecondStage1StageBias12 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=4e-6 W=276e-6
mSimpleFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=12e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=25e-6
mSimpleFirstStageLoad15 FirstStageYout1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=327e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=491e-6
mSimpleFirstStageLoad17 outFirstStage inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=327e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11e-12
.EOM two_stage_single_output_op_amp_195_8

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 3.29901 mW
** Area: 6277 (mu_m)^2
** Transit frequency: 4.55301 MHz
** Transit frequency with error factor: 4.53141 MHz
** Slew rate: 4.29059 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.82001 V
** VoutMin: 0.780001 V
** VcmMax: 5.24001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 3.82581e+07 muA
** DiodeTransistorNmos: 1.37699e+08 muA
** DiodeTransistorNmos: 1.377e+08 muA
** NormalTransistorNmos: 1.37699e+08 muA
** NormalTransistorNmos: 1.377e+08 muA
** NormalTransistorPmos: -1.61506e+08 muA
** NormalTransistorPmos: -1.61506e+08 muA
** NormalTransistorNmos: 4.76151e+07 muA
** NormalTransistorNmos: 4.76141e+07 muA
** NormalTransistorNmos: 2.38081e+07 muA
** NormalTransistorNmos: 2.38081e+07 muA
** NormalTransistorNmos: 2.88581e+08 muA
** NormalTransistorNmos: 2.8858e+08 muA
** NormalTransistorPmos: -2.8858e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -3.82589e+07 muA


** Expected Voltages: 
** ibias: 1.11701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 4.26901  V
** out: 2.5  V
** outFirstStage: 4.25401  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.11601  V
** innerStageBias: 0.557001  V
** innerTransistorStack2Load1: 1.11601  V
** out1: 2.26101  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.489001  V


.END