** Name: two_stage_single_output_op_amp_75_7

.MACRO two_stage_single_output_op_amp_75_7 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=45e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=40e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=13e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=584e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=59e-6
m8 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
m9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=40e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=32e-6
m11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=32e-6
m12 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=56e-6
m13 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=421e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=316e-6
m15 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=80e-6
m16 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=28e-6
m17 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=80e-6
m18 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=41e-6
m19 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=41e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_75_7

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 5.69201 mW
** Area: 8674 (mu_m)^2
** Transit frequency: 3.30601 MHz
** Transit frequency with error factor: 3.30563 MHz
** Slew rate: 3.58089 V/mu_s
** Phase margin: 65.8902°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 0.310001 V
** VcmMax: 5.15001 V
** VcmMin: 1.45001 V


** Expected Currents: 
** NormalTransistorPmos: -2.5096e+08 muA
** NormalTransistorPmos: -1.63609e+07 muA
** NormalTransistorPmos: -1.62449e+07 muA
** NormalTransistorPmos: -2.44399e+07 muA
** NormalTransistorPmos: -1.62449e+07 muA
** NormalTransistorPmos: -2.44399e+07 muA
** DiodeTransistorNmos: 1.62441e+07 muA
** NormalTransistorNmos: 1.62441e+07 muA
** NormalTransistorNmos: 1.62441e+07 muA
** NormalTransistorNmos: 1.63871e+07 muA
** NormalTransistorNmos: 1.63861e+07 muA
** NormalTransistorNmos: 8.19401e+06 muA
** NormalTransistorNmos: 8.19401e+06 muA
** NormalTransistorNmos: 8.02119e+08 muA
** NormalTransistorPmos: -8.02118e+08 muA
** DiodeTransistorNmos: 2.50961e+08 muA
** DiodeTransistorNmos: 1.63601e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.08101  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.17901  V
** outVoltageBiasXXnXX2: 0.716001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.520001  V
** innerTransistorStack2Load2: 0.525001  V
** out1: 0.588001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.92101  V


.END