** Name: symmetrical_op_amp25

.MACRO symmetrical_op_amp25 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mSecondStage1StageBias3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
mSymmetricalFirstStageLoad4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=460e-6
mMainBias5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=8e-6
mSymmetricalFirstStageLoad6 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=460e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=147e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias9 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=147e-6
mMainBias10 inOutputTransconductanceComplementarySecondStage ibias sourceNmos sourceNmos nmos4 L=4e-6 W=16e-6
mSymmetricalFirstStageTransconductor11 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias12 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=3e-6 W=161e-6
mMainBias13 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
mSecondStage1StageBias14 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=159e-6
mSymmetricalFirstStageTransconductor15 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=598e-6
mMainBias18 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=48e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor19 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=3e-6 W=174e-6
mSecondStage1Transconductor20 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=174e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp25

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 6.13601 mW
** Area: 7978 (mu_m)^2
** Transit frequency: 9.51101 MHz
** Transit frequency with error factor: 9.51107 MHz
** Slew rate: 32.9403 V/mu_s
** Phase margin: 76.7764°
** CMRR: 135 dB
** negPSRR: 37 dB
** posPSRR: 32 dB
** VoutMax: 4.26001 V
** VoutMin: 0.550001 V
** VcmMax: 4.67001 V
** VcmMin: 1.15001 V


** Expected Currents: 
** NormalTransistorNmos: 5.75101e+06 muA
** NormalTransistorNmos: 1.34081e+07 muA
** NormalTransistorPmos: -3.40519e+07 muA
** DiodeTransistorPmos: -2.5141e+08 muA
** DiodeTransistorPmos: -2.5141e+08 muA
** NormalTransistorNmos: 5.0282e+08 muA
** NormalTransistorNmos: 2.51411e+08 muA
** NormalTransistorNmos: 2.51411e+08 muA
** NormalTransistorNmos: 3.30573e+08 muA
** NormalTransistorNmos: 3.30572e+08 muA
** NormalTransistorPmos: -3.30572e+08 muA
** NormalTransistorPmos: -3.30571e+08 muA
** NormalTransistorNmos: 3.30573e+08 muA
** NormalTransistorNmos: 3.30572e+08 muA
** NormalTransistorPmos: -3.30572e+08 muA
** NormalTransistorPmos: -3.30571e+08 muA
** DiodeTransistorNmos: 3.40511e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.75199e+06 muA
** DiodeTransistorPmos: -1.34089e+07 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.957001  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 4.26101  V
** innerComplementarySecondStage: 0.686001  V
** inputVoltageBiasXXpXX0: 3.90701  V
** out: 2.5  V
** outFirstStage: 4.26101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.54801  V
** innerStageBias: 0.281001  V
** innerTransconductance: 4.81201  V
** inner: 0.281001  V
** inner: 4.81201  V


.END