.suckt  two_stage_single_output_op_amp_131_4 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias2 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
mMainBias3 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
mSimpleFirstStageLoad4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad5 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad7 FirstStageYinnerSourceLoad1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageLoad8 outFirstStage outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor10 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1Transconductor12 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
mSecondStage1Transconductor13 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias14 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mSecondStage1StageBias15 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos
mSecondStage1StageBias16 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias17 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias18 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mMainBias19 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_131_4

