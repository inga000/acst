.suckt  symmetrical_op_amp95 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_MainBias_1 inOutputStageBiasComplementarySecondStage outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m_Symmetrical_MainBias_3 out2FirstStage ibias sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_4 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m_Symmetrical_FirstStage_Load_5 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Load_6 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m_Symmetrical_FirstStage_Load_7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_StageBias_8 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Transconductor_9 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_Symmetrical_FirstStage_Transconductor_10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_Transconductor_11 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_Symmetrical_SecondStage1_Transconductor_12 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_StageBias_13 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m_Symmetrical_SecondStage1_StageBias_14 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_15 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_16 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_17 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_19 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_20 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_21 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_MainBias_22 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp95

