** Name: two_stage_single_output_op_amp_32_7

.MACRO two_stage_single_output_op_amp_32_7 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=22e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
m4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=5e-6 W=151e-6
m5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=101e-6
m6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=38e-6
m7 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=11e-6
m8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=22e-6
m9 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=9e-6
m10 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=506e-6
m11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=38e-6
m12 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=5e-6 W=151e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=373e-6
m14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=10e-6 W=91e-6
m15 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=442e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.30001e-12
.EOM two_stage_single_output_op_amp_32_7

** Expected Performance Values: 
** Gain: 88 dB
** Power consumption: 3.62701 mW
** Area: 10702 (mu_m)^2
** Transit frequency: 3.52501 MHz
** Transit frequency with error factor: 3.52219 MHz
** Slew rate: 3.86406 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** negPSRR: 96 dB
** posPSRR: 93 dB
** VoutMax: 4.25 V
** VoutMin: 0.210001 V
** VcmMax: 4.42001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorNmos: 1.12661e+07 muA
** NormalTransistorPmos: -4.83919e+07 muA
** NormalTransistorPmos: -1.22419e+07 muA
** NormalTransistorPmos: -1.22419e+07 muA
** DiodeTransistorPmos: -1.22419e+07 muA
** NormalTransistorNmos: 2.44811e+07 muA
** DiodeTransistorNmos: 2.44801e+07 muA
** NormalTransistorNmos: 1.22411e+07 muA
** NormalTransistorNmos: 1.22411e+07 muA
** NormalTransistorNmos: 6.31203e+08 muA
** NormalTransistorPmos: -6.31202e+08 muA
** DiodeTransistorNmos: 4.83911e+07 muA
** NormalTransistorNmos: 4.83911e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.12669e+07 muA


** Expected Voltages: 
** ibias: 0.615001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.22801  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.13401  V
** outSourceVoltageBiasXXnXX1: 0.567001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.28601  V
** out1: 3.44901  V
** sourceTransconductance: 1.92001  V
** inner: 0.567001  V


.END