.suckt  symmetrical_op_amp17 ibias in1 in2 out sourceNmos sourcePmos
mSymmetricalFirstStageLoad1 outFirstStage outFirstStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad2 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageStageBias3 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSymmetricalFirstStageTransconductor4 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSymmetricalFirstStageTransconductor5 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1StageBias6 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
mSecondStage1StageBias7 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStage1Transconductor8 out outFirstStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias9 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos
mSecondStageWithVoltageBiasAsStageBiasStageBias10 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mMainBias12 ibias ibias sourceNmos sourceNmos nmos
.end symmetrical_op_amp17

