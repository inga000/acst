** Name: two_stage_single_output_op_amp_43_9

.MACRO two_stage_single_output_op_amp_43_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=17e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=8e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=84e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=23e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=9e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=8e-6 W=142e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=56e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=56e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
mSecondStage1StageBias11 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=84e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=91e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=91e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=8e-6 W=252e-6
mMainBias16 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=155e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=129e-6
mFoldedCascodeFirstStageLoad18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=9e-6
mMainBias19 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=8e-6 W=562e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.80001e-12
.EOM two_stage_single_output_op_amp_43_9

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 2.76501 mW
** Area: 13433 (mu_m)^2
** Transit frequency: 2.51801 MHz
** Transit frequency with error factor: 2.51211 MHz
** Slew rate: 3.6987 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 1.79001 V
** VcmMax: 4.03001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -4.00199e+07 muA
** NormalTransistorPmos: -1.09519e+07 muA
** NormalTransistorNmos: 1.77771e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** NormalTransistorNmos: 1.77771e+07 muA
** NormalTransistorNmos: 2.66651e+07 muA
** DiodeTransistorPmos: -1.77779e+07 muA
** NormalTransistorPmos: -1.77779e+07 muA
** NormalTransistorPmos: -1.77789e+07 muA
** NormalTransistorPmos: -8.88899e+06 muA
** NormalTransistorPmos: -8.88899e+06 muA
** NormalTransistorNmos: 4.28684e+08 muA
** DiodeTransistorNmos: 4.28683e+08 muA
** NormalTransistorPmos: -4.28683e+08 muA
** DiodeTransistorNmos: 4.00191e+07 muA
** NormalTransistorNmos: 4.00191e+07 muA
** DiodeTransistorNmos: 1.09511e+07 muA
** DiodeTransistorNmos: 1.09521e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.13401  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 2.19201  V
** outSourceVoltageBiasXXnXX1: 1.09601  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.68901  V
** sourceGCC1: 0.528001  V
** sourceGCC2: 0.528001  V
** sourceTransconductance: 3.29701  V
** inner: 1.09601  V


.END