.suckt  two_stage_fully_differential_op_amp_56_11 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m3 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m5 outFeedback outFeedback sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m7 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m8 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m9 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m14 out1FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m15 FirstStageYinnerTransistorStack1Load1 outFeedback sourcePmos sourcePmos pmos
m16 out2FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m17 FirstStageYinnerTransistorStack2Load1 outFeedback sourcePmos sourcePmos pmos
m18 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m19 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m20 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m21 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m22 out1 ibias SecondStage1YinnerStageBias SecondStage1YinnerStageBias nmos
m23 SecondStage1YinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m24 out1 outVoltageBiasXXpXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
m25 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m26 out2 ibias SecondStage2YinnerStageBias SecondStage2YinnerStageBias nmos
m27 SecondStage2YinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m28 out2 outVoltageBiasXXpXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
m29 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
m30 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m31 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m32 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m33 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m34 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m35 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_56_11

