** Name: two_stage_single_output_op_amp_60_1

.MACRO two_stage_single_output_op_amp_60_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=17e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=16e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=175e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=16e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=28e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=116e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=116e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=65e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=28e-6
mMainBias12 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=100e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=64e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=64e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=175e-6
mMainBias18 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=16e-6
mSecondStage1StageBias19 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=530e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=9e-6 W=231e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_60_1

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 4.95401 mW
** Area: 10055 (mu_m)^2
** Transit frequency: 4.47001 MHz
** Transit frequency with error factor: 4.4702 MHz
** Slew rate: 4.60383 V/mu_s
** Phase margin: 63.5984°
** CMRR: 141 dB
** VoutMax: 4.31001 V
** VoutMin: 0.570001 V
** VcmMax: 3.37001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.94901e+06 muA
** NormalTransistorNmos: 2.73401e+07 muA
** NormalTransistorNmos: 2.09531e+07 muA
** NormalTransistorNmos: 3.16681e+07 muA
** NormalTransistorNmos: 2.09531e+07 muA
** NormalTransistorNmos: 3.16681e+07 muA
** NormalTransistorPmos: -2.09539e+07 muA
** NormalTransistorPmos: -2.09539e+07 muA
** DiodeTransistorPmos: -2.09539e+07 muA
** NormalTransistorPmos: -2.14329e+07 muA
** DiodeTransistorPmos: -2.14339e+07 muA
** NormalTransistorPmos: -1.07159e+07 muA
** NormalTransistorPmos: -1.07159e+07 muA
** NormalTransistorNmos: 8.881e+08 muA
** NormalTransistorPmos: -8.88099e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.94999e+06 muA
** NormalTransistorPmos: -1.95099e+06 muA
** DiodeTransistorPmos: -2.73409e+07 muA


** Expected Voltages: 
** ibias: 1.18101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.976001  V
** outInputVoltageBiasXXpXX1: 3.54001  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outSourceVoltageBiasXXpXX1: 4.27001  V
** outVoltageBiasXXpXX2: 3.74801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.25  V
** out1: 3.47201  V
** sourceGCC1: 0.526001  V
** sourceGCC2: 0.526001  V
** sourceTransconductance: 3.23101  V
** inner: 4.26901  V


.END