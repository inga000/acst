** Name: two_stage_single_output_op_amp_62_1

.MACRO two_stage_single_output_op_amp_62_1 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=13e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
m3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=6e-6 W=14e-6
m5 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
m6 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=22e-6
m7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
m8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=37e-6
m9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=147e-6
m10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=147e-6
m11 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=62e-6
m12 inputVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=50e-6
m13 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=156e-6
m14 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=37e-6
m15 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=102e-6
m16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=132e-6
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=132e-6
m19 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=21e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
m21 out inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=2e-6 W=366e-6
m22 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=375e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 5.40001e-12
.EOM two_stage_single_output_op_amp_62_1

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 4.47301 mW
** Area: 9129 (mu_m)^2
** Transit frequency: 4.62101 MHz
** Transit frequency with error factor: 4.62065 MHz
** Slew rate: 6.79531 V/mu_s
** Phase margin: 60.1606°
** CMRR: 137 dB
** VoutMax: 4.54001 V
** VoutMin: 0.560001 V
** VcmMax: 3 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.91141e+07 muA
** NormalTransistorNmos: 2.36901e+07 muA
** NormalTransistorNmos: 1.91791e+07 muA
** NormalTransistorNmos: 3.72281e+07 muA
** NormalTransistorNmos: 5.59961e+07 muA
** NormalTransistorNmos: 3.72281e+07 muA
** NormalTransistorNmos: 5.59961e+07 muA
** DiodeTransistorPmos: -3.72289e+07 muA
** NormalTransistorPmos: -3.72289e+07 muA
** NormalTransistorPmos: -3.72289e+07 muA
** NormalTransistorPmos: -3.75389e+07 muA
** DiodeTransistorPmos: -3.75399e+07 muA
** NormalTransistorPmos: -1.87689e+07 muA
** NormalTransistorPmos: -1.87689e+07 muA
** NormalTransistorNmos: 6.90711e+08 muA
** NormalTransistorPmos: -6.9071e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.91149e+07 muA
** NormalTransistorPmos: -3.91159e+07 muA
** DiodeTransistorPmos: -2.36909e+07 muA
** DiodeTransistorPmos: -1.91799e+07 muA


** Expected Voltages: 
** ibias: 1.17301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.68601  V
** inputVoltageBiasXXpXX3: 3.97501  V
** out: 2.5  V
** outFirstStage: 0.968001  V
** outInputVoltageBiasXXpXX1: 3.23801  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.11901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.43201  V
** out1: 4.18801  V
** sourceGCC1: 0.523001  V
** sourceGCC2: 0.523001  V
** sourceTransconductance: 3.29901  V
** inner: 4.11601  V


.END