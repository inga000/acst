.suckt  complementary_op_amp34 ibias in1 in2 out sourceNmos sourcePmos
m_Complementary_MainBias_1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_MainBias_2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_3 FirstStageYinnerOutputLoadNmos outInputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m_Complementary_FirstStage_Load_4 FirstStageYinnerTransistorStack1LoadPmos outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_5 out outInputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m_Complementary_FirstStage_Load_6 FirstStageYinnerTransistorStack2LoadPmos outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_7 FirstStageYinnerOutputLoadNmos FirstStageYinnerOutputLoadNmos FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m_Complementary_FirstStage_Load_8 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_9 out FirstStageYinnerOutputLoadNmos FirstStageYinnerSourceLoadNmos FirstStageYinnerSourceLoadNmos nmos
m_Complementary_FirstStage_Load_10 FirstStageYinnerSourceLoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_11 FirstStageYsourceTransconductanceNmos ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_Complementary_FirstStage_StageBias_12 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_13 FirstStageYsourceTransconductancePmos outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_Complementary_FirstStage_StageBias_14 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Transconductor_15 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_16 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_17 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m_Complementary_FirstStage_Transconductor_18 FirstStageYinnerSourceLoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c_Complementary_Load_Capacitor_1 out sourceNmos 
m_Complementary_MainBias_19 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_Complementary_MainBias_20 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_MainBias_21 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_Complementary_MainBias_22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_MainBias_23 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m_Complementary_MainBias_24 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end complementary_op_amp34

