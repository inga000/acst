** Name: two_stage_single_output_op_amp_74_8

.MACRO two_stage_single_output_op_amp_74_8 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=36e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=29e-6
mMainBias3 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=6e-6 W=17e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=26e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=24e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=9e-6 W=36e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=28e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=28e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=26e-6
mSecondStage1StageBias12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=370e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=29e-6
mSecondStage1StageBias14 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=6e-6 W=166e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=174e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=75e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=75e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=536e-6
mFoldedCascodeFirstStageLoad20 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=174e-6
mMainBias21 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=60e-6
mMainBias22 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=100e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6e-12
.EOM two_stage_single_output_op_amp_74_8

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 5.38301 mW
** Area: 10255 (mu_m)^2
** Transit frequency: 3.46501 MHz
** Transit frequency with error factor: 3.46545 MHz
** Slew rate: 3.88913 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 1.44001 V
** VcmMax: 5.12001 V
** VcmMin: 1.43001 V


** Expected Currents: 
** NormalTransistorPmos: -2.86569e+07 muA
** NormalTransistorPmos: -4.81179e+07 muA
** NormalTransistorPmos: -2.35549e+07 muA
** NormalTransistorPmos: -3.63969e+07 muA
** NormalTransistorPmos: -2.35549e+07 muA
** NormalTransistorPmos: -3.63969e+07 muA
** NormalTransistorNmos: 2.35541e+07 muA
** NormalTransistorNmos: 2.35541e+07 muA
** DiodeTransistorNmos: 2.35541e+07 muA
** NormalTransistorNmos: 2.56811e+07 muA
** DiodeTransistorNmos: 2.56801e+07 muA
** NormalTransistorNmos: 1.28411e+07 muA
** NormalTransistorNmos: 1.28411e+07 muA
** NormalTransistorNmos: 9.07037e+08 muA
** NormalTransistorNmos: 9.07036e+08 muA
** NormalTransistorPmos: -9.07036e+08 muA
** DiodeTransistorNmos: 2.86561e+07 muA
** NormalTransistorNmos: 2.86551e+07 muA
** DiodeTransistorNmos: 4.81171e+07 muA
** DiodeTransistorNmos: 4.81161e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.24001  V
** outInputVoltageBiasXXnXX2: 1.67101  V
** outSourceVoltageBiasXXnXX1: 0.620001  V
** outSourceVoltageBiasXXnXX2: 0.820001  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.668001  V
** out1: 1.22501  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.90001  V
** innerStageBias: 0.641001  V
** inner: 0.618001  V


.END