** Name: two_stage_single_output_op_amp_3_2

.MACRO two_stage_single_output_op_amp_3_2 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=101e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
m4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=4e-6 W=101e-6
m5 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=108e-6
m6 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=3e-6 W=118e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=50e-6
m8 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=38e-6
m9 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=181e-6
m10 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=34e-6
m11 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=392e-6
m12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=38e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_3_2

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 1.71201 mW
** Area: 2666 (mu_m)^2
** Transit frequency: 4.49901 MHz
** Transit frequency with error factor: 4.48618 MHz
** Slew rate: 8.44558 V/mu_s
** Phase margin: 65.8902°
** CMRR: 92 dB
** negPSRR: 90 dB
** posPSRR: 96 dB
** VoutMax: 4.83001 V
** VoutMin: 0.400001 V
** VcmMax: 3.51001 V
** VcmMin: 0.180001 V


** Expected Currents: 
** NormalTransistorPmos: -1.81499e+07 muA
** DiodeTransistorNmos: 4.82271e+07 muA
** NormalTransistorNmos: 4.82271e+07 muA
** NormalTransistorNmos: 4.82271e+07 muA
** NormalTransistorPmos: -9.64569e+07 muA
** NormalTransistorPmos: -4.82279e+07 muA
** NormalTransistorPmos: -4.82279e+07 muA
** NormalTransistorNmos: 2.07779e+08 muA
** NormalTransistorNmos: 2.07778e+08 muA
** NormalTransistorPmos: -2.07778e+08 muA
** DiodeTransistorNmos: 1.81491e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.804001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack2Load1: 0.214001  V
** sourceTransconductance: 3.81401  V
** innerTransconductance: 0.150001  V


.END