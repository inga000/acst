.suckt  symmetrical_op_amp153 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_MainBias_1 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_2 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m_Symmetrical_FirstStage_Load_3 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Load_4 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m_Symmetrical_FirstStage_Load_5 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_StageBias_6 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_Symmetrical_FirstStage_StageBias_7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Transconductor_8 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_Symmetrical_FirstStage_Transconductor_9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_Transconductor_10 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_Symmetrical_SecondStage1_Transconductor_11 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_StageBias_12 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos
m_Symmetrical_SecondStage1_StageBias_13 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_14 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_15 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_17 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_18 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_Symmetrical_MainBias_19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end symmetrical_op_amp153

