.suckt  symmetrical_op_amp13 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_MainBias_1 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_2 outFirstStage outFirstStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Load_3 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_StageBias_4 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Transconductor_5 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_Symmetrical_FirstStage_Transconductor_6 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_Transconductor_7 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_Symmetrical_SecondStage1_Transconductor_8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_StageBias_9 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos
m_Symmetrical_SecondStage1_StageBias_10 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_11 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_12 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_13 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_StageBias_14 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_15 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp13

