.suckt  one_stage_fully_differential_op_amp17 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
m1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m3 outFeedback outFeedback sourcePmos sourcePmos pmos
m4 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m5 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m6 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m7 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m8 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m9 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m10 out1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m11 FirstStageYsourceGCC1 outFeedback sourcePmos sourcePmos pmos
m12 out2 inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m13 FirstStageYsourceGCC2 outFeedback sourcePmos sourcePmos pmos
m14 out1 ibias sourceNmos sourceNmos nmos
m15 out2 ibias sourceNmos sourceNmos nmos
m16 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out1 sourceNmos 
c2 out2 sourceNmos 
m19 ibias ibias sourceNmos sourceNmos nmos
m20 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end one_stage_fully_differential_op_amp17

