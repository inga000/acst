** Name: two_stage_single_output_op_amp_16_1

.MACRO two_stage_single_output_op_amp_16_1 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
m2 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=58e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=21e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=14e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=137e-6
m6 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=219e-6
m7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=58e-6
m8 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=10e-6
m9 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=6e-6
m10 out ibias sourcePmos sourcePmos pmos4 L=6e-6 W=288e-6
m11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=72e-6
m12 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=72e-6
m13 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=137e-6
m14 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=14e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_16_1

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 0.962001 mW
** Area: 5747 (mu_m)^2
** Transit frequency: 3.82001 MHz
** Transit frequency with error factor: 3.81169 MHz
** Slew rate: 5.65174 V/mu_s
** Phase margin: 64.1713°
** CMRR: 97 dB
** negPSRR: 98 dB
** posPSRR: 210 dB
** VoutMax: 4.60001 V
** VoutMin: 0.150001 V
** VcmMax: 3.19001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 2.86401e+06 muA
** NormalTransistorPmos: -2.89499e+06 muA
** DiodeTransistorNmos: 1.38091e+07 muA
** NormalTransistorNmos: 1.38091e+07 muA
** NormalTransistorPmos: -2.76189e+07 muA
** DiodeTransistorPmos: -2.76199e+07 muA
** NormalTransistorPmos: -1.38099e+07 muA
** NormalTransistorPmos: -1.38099e+07 muA
** NormalTransistorNmos: 1.39052e+08 muA
** NormalTransistorPmos: -1.39051e+08 muA
** DiodeTransistorNmos: 2.89401e+06 muA
** DiodeTransistorPmos: -2.86499e+06 muA
** NormalTransistorPmos: -2.86599e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.03501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.589001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.44601  V
** outSourceVoltageBiasXXpXX1: 4.22301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceTransconductance: 3.31701  V
** inner: 4.22301  V


.END