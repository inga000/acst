** Name: two_stage_single_output_op_amp_43_7

.MACRO two_stage_single_output_op_amp_43_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=60e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=115e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=74e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=74e-6
mSecondStage1StageBias8 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mFoldedCascodeFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=115e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=279e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=279e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=5e-6 W=600e-6
mMainBias13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=159e-6
mSecondStage1Transconductor14 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=411e-6
mFoldedCascodeFirstStageLoad15 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=30e-6
mMainBias16 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=125e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 17.6001e-12
.EOM two_stage_single_output_op_amp_43_7

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 7.52101 mW
** Area: 8799 (mu_m)^2
** Transit frequency: 5.25701 MHz
** Transit frequency with error factor: 5.25156 MHz
** Slew rate: 5.102 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.60001 V
** VoutMin: 0.150001 V
** VcmMax: 4.04001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.70289e+07 muA
** NormalTransistorPmos: -2.09519e+07 muA
** NormalTransistorNmos: 8.99431e+07 muA
** NormalTransistorNmos: 1.40944e+08 muA
** NormalTransistorNmos: 8.99431e+07 muA
** NormalTransistorNmos: 1.40944e+08 muA
** DiodeTransistorPmos: -8.99439e+07 muA
** NormalTransistorPmos: -8.99439e+07 muA
** NormalTransistorPmos: -1.01996e+08 muA
** NormalTransistorPmos: -5.09989e+07 muA
** NormalTransistorPmos: -5.09989e+07 muA
** NormalTransistorNmos: 1.15432e+09 muA
** NormalTransistorPmos: -1.15431e+09 muA
** DiodeTransistorNmos: 2.70281e+07 muA
** DiodeTransistorNmos: 2.09511e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.969001  V
** out: 2.5  V
** outFirstStage: 4.03801  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.02501  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.23901  V


.END