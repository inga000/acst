** Name: two_stage_single_output_op_amp_9_8

.MACRO two_stage_single_output_op_amp_9_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=11e-6
m3 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=11e-6
m4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=43e-6
m5 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=126e-6
m6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=14e-6
m7 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=14e-6
m9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
m10 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=310e-6
m11 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=202e-6
m12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=2e-6 W=11e-6
m13 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=220e-6
m14 FirstStageYout1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=7e-6 W=43e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_9_8

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 3.61201 mW
** Area: 3883 (mu_m)^2
** Transit frequency: 3.02901 MHz
** Transit frequency with error factor: 3.02454 MHz
** Slew rate: 6.19712 V/mu_s
** Phase margin: 62.4525°
** CMRR: 95 dB
** negPSRR: 95 dB
** posPSRR: 87 dB
** VoutMax: 4.25 V
** VoutMin: 0.420001 V
** VcmMax: 4.11001 V
** VcmMin: 0.930001 V


** Expected Currents: 
** NormalTransistorNmos: 8.21501e+06 muA
** NormalTransistorPmos: -1.63552e+08 muA
** NormalTransistorPmos: -1.39649e+07 muA
** NormalTransistorPmos: -1.39649e+07 muA
** DiodeTransistorPmos: -1.39649e+07 muA
** NormalTransistorNmos: 2.79291e+07 muA
** NormalTransistorNmos: 1.39641e+07 muA
** NormalTransistorNmos: 1.39641e+07 muA
** NormalTransistorNmos: 5.12747e+08 muA
** NormalTransistorNmos: 5.12746e+08 muA
** NormalTransistorPmos: -5.12746e+08 muA
** DiodeTransistorNmos: 1.63553e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.21599e+06 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 0.822001  V
** outVoltageBiasXXpXX0: 3.93401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.08001  V
** out1: 3.14001  V
** sourceTransconductance: 1.76801  V
** innerStageBias: 0.198001  V


.END