.suckt  complementary_op_amp3 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 FirstStageYinnerOutputLoadPmos FirstStageYinnerOutputLoadPmos FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m3 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m4 out FirstStageYinnerOutputLoadPmos FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos pmos
m5 FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m6 FirstStageYinnerOutputLoadPmos FirstStageYinnerOutputLoadPmos FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m7 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m8 out FirstStageYinnerOutputLoadPmos FirstStageYinnerSourceLoadNmos FirstStageYinnerSourceLoadNmos nmos
m9 FirstStageYinnerSourceLoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m10 FirstStageYsourceTransconductanceNmos inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m11 FirstStageYsourceTransconductancePmos ibias sourcePmos sourcePmos pmos
m12 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m13 FirstStageYinnerSourceLoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m14 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m15 FirstStageYinnerSourceLoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c1 out sourceNmos 
m16 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m17 ibias ibias sourcePmos sourcePmos pmos
.end complementary_op_amp3

