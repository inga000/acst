** Name: two_stage_single_output_op_amp_10_10

.MACRO two_stage_single_output_op_amp_10_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
m2 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=43e-6
m3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=320e-6
m4 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=16e-6
m5 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=491e-6
m6 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=241e-6
m7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=16e-6
m8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=84e-6
m9 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=64e-6
m10 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=526e-6
m11 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=320e-6
m12 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=495e-6
Capacitor1 outFirstStage out 12.7001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_10_10

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 3.71501 mW
** Area: 8415 (mu_m)^2
** Transit frequency: 2.82301 MHz
** Transit frequency with error factor: 2.81953 MHz
** Slew rate: 5.91017 V/mu_s
** Phase margin: 60.1606°
** CMRR: 102 dB
** negPSRR: 112 dB
** posPSRR: 95 dB
** VoutMax: 4.25 V
** VoutMin: 0.180001 V
** VcmMax: 4.42001 V
** VcmMin: 0.920001 V


** Expected Currents: 
** NormalTransistorNmos: 2.18298e+08 muA
** DiodeTransistorPmos: -3.75969e+07 muA
** NormalTransistorPmos: -3.75969e+07 muA
** NormalTransistorPmos: -3.75969e+07 muA
** NormalTransistorNmos: 7.51921e+07 muA
** NormalTransistorNmos: 3.75961e+07 muA
** NormalTransistorNmos: 3.75961e+07 muA
** NormalTransistorNmos: 4.39515e+08 muA
** NormalTransistorPmos: -4.39514e+08 muA
** NormalTransistorPmos: -4.39515e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.18297e+08 muA


** Expected Voltages: 
** ibias: 0.584001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.99101  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.50601  V
** out1: 4.27401  V
** sourceTransconductance: 1.76101  V
** innerTransconductance: 4.55501  V


.END