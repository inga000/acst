** Name: symmetrical_op_amp36

.MACRO symmetrical_op_amp36 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=8e-6 W=129e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=129e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=54e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=7e-6 W=57e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=197e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=8e-6 W=197e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=2e-6 W=18e-6
mSecondStage1Transconductor11 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=18e-6
mSymmetricalFirstStageStageBias12 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=61e-6
mSymmetricalFirstStageStageBias13 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=31e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=54e-6
mMainBias15 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=46e-6
mSymmetricalFirstStageTransconductor16 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=106e-6
mSecondStage1StageBias17 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=7e-6 W=531e-6
mSymmetricalFirstStageTransconductor18 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=106e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp36

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 1.11101 mW
** Area: 10968 (mu_m)^2
** Transit frequency: 3.37201 MHz
** Transit frequency with error factor: 3.37247 MHz
** Slew rate: 4.65737 V/mu_s
** Phase margin: 60.1606°
** CMRR: 149 dB
** negPSRR: 47 dB
** posPSRR: 54 dB
** VoutMax: 3.66001 V
** VoutMin: 0.400001 V
** VcmMax: 3.08001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorPmos: -4.66379e+07 muA
** DiodeTransistorNmos: 3.09231e+07 muA
** DiodeTransistorNmos: 3.09231e+07 muA
** NormalTransistorPmos: -6.18469e+07 muA
** NormalTransistorPmos: -6.18459e+07 muA
** NormalTransistorPmos: -3.09239e+07 muA
** NormalTransistorPmos: -3.09239e+07 muA
** NormalTransistorNmos: 4.69011e+07 muA
** NormalTransistorNmos: 4.69021e+07 muA
** NormalTransistorPmos: -4.69019e+07 muA
** NormalTransistorPmos: -4.69029e+07 muA
** DiodeTransistorPmos: -4.69039e+07 muA
** DiodeTransistorPmos: -4.69049e+07 muA
** NormalTransistorNmos: 4.69031e+07 muA
** NormalTransistorNmos: 4.69021e+07 muA
** DiodeTransistorNmos: 4.66371e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.802001  V
** inSourceStageBiasComplementarySecondStage: 3.85001  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 2.71601  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.29501  V
** sourceTransconductance: 3.28501  V
** innerStageBias: 3.46601  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END