.suckt  two_stage_single_output_op_amp_111_4 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_3 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_4 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m_SingleOutput_FirstStage_Load_5 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m_SingleOutput_FirstStage_Load_6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m_SingleOutput_FirstStage_Load_7 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_8 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m_SingleOutput_FirstStage_Load_9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_StageBias_10 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m_SingleOutput_FirstStage_StageBias_11 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Transconductor_12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m_SingleOutput_FirstStage_Transconductor_13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_Transconductor_14 out outVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_SingleOutput_SecondStage1_Transconductor_15 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_16 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m_SingleOutput_SecondStage1_StageBias_17 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_18 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_19 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_20 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
m_SingleOutput_MainBias_21 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m_SingleOutput_MainBias_22 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_111_4

