** Name: two_stage_single_output_op_amp_47_5

.MACRO two_stage_single_output_op_amp_47_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=10e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=18e-6
mMainBias4 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=10e-6 W=283e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=19e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=205e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=15e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mMainBias10 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=26e-6
mMainBias11 inputVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=17e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=177e-6
mFoldedCascodeFirstStageLoad13 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=15e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=45e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=7e-6 W=160e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=75e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=8e-6 W=75e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=149e-6
mFoldedCascodeFirstStageTransconductor19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=149e-6
mFoldedCascodeFirstStageStageBias20 FirstStageYsourceTransconductance inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=10e-6 W=331e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=205e-6
mFoldedCascodeFirstStageLoad23 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=160e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_47_5

** Expected Performance Values: 
** Gain: 132 dB
** Power consumption: 3.14301 mW
** Area: 14496 (mu_m)^2
** Transit frequency: 4.25101 MHz
** Transit frequency with error factor: 4.25109 MHz
** Slew rate: 4.15032 V/mu_s
** Phase margin: 60.7336°
** CMRR: 140 dB
** VoutMax: 3.41001 V
** VoutMin: 0.510001 V
** VcmMax: 4.10001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.41441e+07 muA
** NormalTransistorNmos: 2.60201e+07 muA
** NormalTransistorNmos: 1.66771e+07 muA
** NormalTransistorNmos: 1.88141e+07 muA
** NormalTransistorNmos: 2.84491e+07 muA
** NormalTransistorNmos: 1.88141e+07 muA
** NormalTransistorNmos: 2.84491e+07 muA
** NormalTransistorPmos: -1.88149e+07 muA
** NormalTransistorPmos: -1.88159e+07 muA
** NormalTransistorPmos: -1.88149e+07 muA
** NormalTransistorPmos: -1.88159e+07 muA
** NormalTransistorPmos: -1.92729e+07 muA
** NormalTransistorPmos: -9.63599e+06 muA
** NormalTransistorPmos: -9.63599e+06 muA
** NormalTransistorNmos: 4.74779e+08 muA
** NormalTransistorPmos: -4.74778e+08 muA
** DiodeTransistorPmos: -4.74779e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -4.41449e+07 muA
** NormalTransistorPmos: -4.41459e+07 muA
** DiodeTransistorPmos: -2.60209e+07 muA
** DiodeTransistorPmos: -1.66779e+07 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.68601  V
** inputVoltageBiasXXpXX3: 4.25501  V
** out: 2.5  V
** outFirstStage: 0.911001  V
** outInputVoltageBiasXXpXX1: 2.85001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 3.92501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.10001  V
** innerTransistorStack1Load2: 4.46401  V
** innerTransistorStack2Load2: 4.46401  V
** sourceGCC1: 0.538001  V
** sourceGCC2: 0.538001  V
** sourceTransconductance: 3.22301  V
** inner: 3.92201  V


.END