** Name: two_stage_single_output_op_amp_47_3

.MACRO two_stage_single_output_op_amp_47_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=9e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=74e-6
mMainBias4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=153e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=14e-6
mFoldedCascodeFirstStageLoad6 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=45e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=45e-6
mMainBias8 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=565e-6
mMainBias9 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=223e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=64e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=14e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerSourceLoad2 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=38e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=101e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=101e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mSecondStage1StageBias18 SecondStageYinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=569e-6
mSecondStage1StageBias19 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=599e-6
mFoldedCascodeFirstStageLoad20 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=38e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_47_3

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 5.67401 mW
** Area: 6273 (mu_m)^2
** Transit frequency: 4.23401 MHz
** Transit frequency with error factor: 4.23432 MHz
** Slew rate: 4.311 V/mu_s
** Phase margin: 61.8795°
** CMRR: 141 dB
** VoutMax: 4.45001 V
** VoutMin: 0.550001 V
** VcmMax: 4.04001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.75676e+08 muA
** NormalTransistorNmos: 1.47368e+08 muA
** NormalTransistorNmos: 1.94511e+07 muA
** NormalTransistorNmos: 2.94301e+07 muA
** NormalTransistorNmos: 1.94511e+07 muA
** NormalTransistorNmos: 2.94301e+07 muA
** NormalTransistorPmos: -1.94519e+07 muA
** NormalTransistorPmos: -1.94529e+07 muA
** NormalTransistorPmos: -1.94519e+07 muA
** NormalTransistorPmos: -1.94529e+07 muA
** NormalTransistorPmos: -1.99609e+07 muA
** NormalTransistorPmos: -9.97999e+06 muA
** NormalTransistorPmos: -9.97999e+06 muA
** NormalTransistorNmos: 5.42836e+08 muA
** NormalTransistorPmos: -5.42835e+08 muA
** NormalTransistorPmos: -5.42836e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.75675e+08 muA
** DiodeTransistorPmos: -1.47367e+08 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** inputVoltageBiasXXpXX2: 4.20501  V
** out: 2.5  V
** outFirstStage: 0.956001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.20201  V
** innerTransistorStack1Load2: 4.48901  V
** innerTransistorStack2Load2: 4.48901  V
** sourceGCC1: 0.533001  V
** sourceGCC2: 0.533001  V
** sourceTransconductance: 3.23001  V
** innerStageBias: 4.56701  V


.END