** Name: two_stage_single_output_op_amp_8_8

.MACRO two_stage_single_output_op_amp_8_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=13e-6
m3 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=36e-6
m4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=8e-6
m5 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=146e-6
m6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=40e-6
m7 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=22e-6
m8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=40e-6
m9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=23e-6
m10 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=564e-6
m11 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=186e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=79e-6
m13 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=8e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 8.80001e-12
.EOM two_stage_single_output_op_amp_8_8

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 5.17901 mW
** Area: 2553 (mu_m)^2
** Transit frequency: 3.77601 MHz
** Transit frequency with error factor: 3.7714 MHz
** Slew rate: 3.66297 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** negPSRR: 138 dB
** posPSRR: 87 dB
** VoutMax: 4.25 V
** VoutMin: 0.540001 V
** VcmMax: 4.09001 V
** VcmMin: 0.740001 V


** Expected Currents: 
** NormalTransistorNmos: 3.14241e+07 muA
** NormalTransistorPmos: -1.60036e+08 muA
** DiodeTransistorPmos: -1.61399e+07 muA
** NormalTransistorPmos: -1.61399e+07 muA
** NormalTransistorNmos: 3.22781e+07 muA
** NormalTransistorNmos: 1.61391e+07 muA
** NormalTransistorNmos: 1.61391e+07 muA
** NormalTransistorNmos: 8.02119e+08 muA
** NormalTransistorNmos: 8.02118e+08 muA
** NormalTransistorPmos: -8.02118e+08 muA
** DiodeTransistorNmos: 1.60037e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.14249e+07 muA


** Expected Voltages: 
** ibias: 0.588001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.947001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 4.125  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.68601  V
** sourceTransconductance: 1.94001  V
** innerStageBias: 0.183001  V


.END