** Name: two_stage_single_output_op_amp_82_7

.MACRO two_stage_single_output_op_amp_82_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=1e-6 W=12e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=34e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=6e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=28e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=12e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=19e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=32e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=32e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=6e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=34e-6
mSecondStage1StageBias13 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=315e-6
mFoldedCascodeFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=12e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=135e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=78e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=78e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=147e-6
mFoldedCascodeFirstStageLoad19 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=135e-6
mMainBias20 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=301e-6
mMainBias21 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=245e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_82_7

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 9.43301 mW
** Area: 5027 (mu_m)^2
** Transit frequency: 5.18401 MHz
** Transit frequency with error factor: 5.18359 MHz
** Slew rate: 6.03242 V/mu_s
** Phase margin: 67.0361°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 0.580001 V
** VcmMax: 5.16001 V
** VcmMin: 1.94001 V


** Expected Currents: 
** NormalTransistorPmos: -1.60411e+08 muA
** NormalTransistorPmos: -1.30567e+08 muA
** NormalTransistorPmos: -2.74139e+07 muA
** NormalTransistorPmos: -4.15679e+07 muA
** NormalTransistorPmos: -2.74139e+07 muA
** NormalTransistorPmos: -4.15679e+07 muA
** DiodeTransistorNmos: 2.74131e+07 muA
** NormalTransistorNmos: 2.74121e+07 muA
** NormalTransistorNmos: 2.74131e+07 muA
** DiodeTransistorNmos: 2.74121e+07 muA
** NormalTransistorNmos: 2.83051e+07 muA
** DiodeTransistorNmos: 2.83041e+07 muA
** NormalTransistorNmos: 1.41531e+07 muA
** NormalTransistorNmos: 1.41531e+07 muA
** NormalTransistorNmos: 1.49256e+09 muA
** NormalTransistorPmos: -1.49255e+09 muA
** DiodeTransistorNmos: 1.60412e+08 muA
** NormalTransistorNmos: 1.60411e+08 muA
** DiodeTransistorNmos: 1.30568e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.75  V
** outSourceVoltageBiasXXnXX1: 0.875  V
** outSourceVoltageBiasXXpXX1: 4.19301  V
** outVoltageBiasXXnXX2: 0.982001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.568001  V
** innerTransistorStack2Load2: 0.569001  V
** out1: 1.13801  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.90301  V
** inner: 0.871001  V


.END