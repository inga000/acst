** Name: one_stage_single_output_op_amp68

.MACRO one_stage_single_output_op_amp68 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=50e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=43e-6
m3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=41e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=301e-6
m5 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=90e-6
m6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=6e-6 W=90e-6
m7 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=39e-6
m8 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=39e-6
m9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=50e-6
m10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=50e-6
m11 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=388e-6
m12 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=90e-6
m13 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=90e-6
m14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=92e-6
m15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=92e-6
m16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=301e-6
m17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=41e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp68

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 1.69001 mW
** Area: 6003 (mu_m)^2
** Transit frequency: 3.92701 MHz
** Transit frequency with error factor: 3.92719 MHz
** Slew rate: 3.70865 V/mu_s
** Phase margin: 89.3815°
** CMRR: 134 dB
** VoutMax: 3.69001 V
** VoutMin: 0.720001 V
** VcmMax: 3.25 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorPmos: -9.52329e+07 muA
** NormalTransistorNmos: 7.42811e+07 muA
** NormalTransistorNmos: 1.11424e+08 muA
** NormalTransistorNmos: 7.42811e+07 muA
** NormalTransistorNmos: 1.11424e+08 muA
** DiodeTransistorPmos: -7.42819e+07 muA
** NormalTransistorPmos: -7.42829e+07 muA
** NormalTransistorPmos: -7.42819e+07 muA
** DiodeTransistorPmos: -7.42829e+07 muA
** NormalTransistorPmos: -7.42869e+07 muA
** DiodeTransistorPmos: -7.42879e+07 muA
** NormalTransistorPmos: -3.71429e+07 muA
** NormalTransistorPmos: -3.71429e+07 muA
** DiodeTransistorNmos: 9.52321e+07 muA
** DiodeTransistorNmos: 9.52311e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.12201  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.567001  V
** outSourceVoltageBiasXXpXX1: 4.20201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.21601  V
** innerTransistorStack2Load2: 4.22101  V
** out1: 3.12801  V
** sourceGCC1: 0.567001  V
** sourceGCC2: 0.567001  V
** sourceTransconductance: 3.21401  V
** inner: 4.19901  V


.END