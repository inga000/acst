.suckt  two_stage_single_output_op_amp_194_10 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
m5 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos
m6 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m7 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourceNmos sourceNmos nmos
m8 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m9 FirstStageYinnerTransistorStack1Load2 ibias sourcePmos sourcePmos pmos
m10 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m11 FirstStageYinnerTransistorStack2Load2 ibias sourcePmos sourcePmos pmos
m12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m13 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m14 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c2 out sourceNmos 
m16 out inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m18 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
m19 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m20 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m21 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m22 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m23 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m24 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_194_10

