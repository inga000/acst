.suckt  two_stage_single_output_op_amp_117_10 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mMainBias2 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mMainBias4 inputVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mTelescopicFirstStageLoad5 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
mTelescopicFirstStageLoad6 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
mTelescopicFirstStageLoad7 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
mTelescopicFirstStageLoad8 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
mTelescopicFirstStageLoad9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos
mTelescopicFirstStageStageBias10 sourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
mTelescopicFirstStageStageBias11 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias14 out ibias sourceNmos sourceNmos nmos
mSecondStage1Transconductor15 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
mMainBias17 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
mMainBias18 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
mMainBias19 ibias ibias sourceNmos sourceNmos nmos
mMainBias20 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mMainBias21 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_117_10

