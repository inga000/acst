** Name: two_stage_single_output_op_amp_9_7

.MACRO two_stage_single_output_op_amp_9_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
mSimpleFirstStageLoad2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSimpleFirstStageTransconductor3 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=12e-6
mSimpleFirstStageStageBias4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias5 out ibias sourceNmos sourceNmos nmos4 L=2e-6 W=305e-6
mSimpleFirstStageTransconductor6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=12e-6
mSimpleFirstStageLoad7 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mSecondStage1Transconductor8 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=102e-6
mSimpleFirstStageLoad9 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=5e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_9_7

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 2.68801 mW
** Area: 1022 (mu_m)^2
** Transit frequency: 2.63501 MHz
** Transit frequency with error factor: 2.63312 MHz
** Slew rate: 3.6473 V/mu_s
** Phase margin: 65.8902°
** CMRR: 97 dB
** negPSRR: 95 dB
** posPSRR: 91 dB
** VoutMax: 4.25 V
** VoutMin: 0.200001 V
** VcmMax: 4.21001 V
** VcmMin: 0.820001 V


** Expected Currents: 
** NormalTransistorPmos: -8.21499e+06 muA
** NormalTransistorPmos: -8.21499e+06 muA
** DiodeTransistorPmos: -8.21499e+06 muA
** NormalTransistorNmos: 1.64291e+07 muA
** NormalTransistorNmos: 8.21401e+06 muA
** NormalTransistorNmos: 8.21401e+06 muA
** NormalTransistorNmos: 5.11202e+08 muA
** NormalTransistorPmos: -5.11201e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load1: 4.23101  V
** out1: 3.23801  V
** sourceTransconductance: 1.87401  V


.END