.suckt  two_stage_fully_differential_op_amp_26_10 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m4 outFeedback outFeedback sourceNmos sourceNmos nmos
m5 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m6 FeedbackStageYinnerStageBias1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m7 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m8 FeedbackStageYinnerStageBias2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m9 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m10 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m11 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m12 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m13 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m14 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m15 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos
m16 FirstStageYinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m17 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m18 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m19 out1 ibias sourceNmos sourceNmos nmos
m20 out1 outVoltageBiasXXpXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
m21 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m22 out2 ibias sourceNmos sourceNmos nmos
m23 out2 outVoltageBiasXXpXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
m24 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
m25 ibias ibias sourceNmos sourceNmos nmos
m26 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m27 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_26_10

