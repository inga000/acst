** Name: symmetrical_op_amp35

.MACRO symmetrical_op_amp35 ibias in1 in2 out sourceNmos sourcePmos
m1 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
m2 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
m3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
m4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=80e-6
m6 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=96e-6
m7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m8 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=32e-6
m9 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=32e-6
m10 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=158e-6
m11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=46e-6
m12 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=46e-6
m13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=39e-6
m14 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=6e-6 W=439e-6
m15 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=147e-6
m16 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=12e-6
m17 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=39e-6
m18 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=182e-6
m19 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=56e-6
m20 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=96e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp35

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 1.42801 mW
** Area: 7665 (mu_m)^2
** Transit frequency: 3.05801 MHz
** Transit frequency with error factor: 3.05838 MHz
** Slew rate: 3.5 V/mu_s
** Phase margin: 69.328°
** CMRR: 142 dB
** negPSRR: 52 dB
** posPSRR: 65 dB
** VoutMax: 4.35001 V
** VoutMin: 0.510001 V
** VcmMax: 3.34001 V
** VcmMin: 0.0700001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00312e+08 muA
** NormalTransistorPmos: -1.85849e+07 muA
** NormalTransistorPmos: -5.45e+07 muA
** DiodeTransistorNmos: 1.12781e+07 muA
** DiodeTransistorNmos: 1.12781e+07 muA
** NormalTransistorPmos: -2.25589e+07 muA
** NormalTransistorPmos: -2.25599e+07 muA
** NormalTransistorPmos: -1.12789e+07 muA
** NormalTransistorPmos: -1.12789e+07 muA
** NormalTransistorNmos: 3.50161e+07 muA
** NormalTransistorNmos: 3.50151e+07 muA
** NormalTransistorPmos: -3.50169e+07 muA
** NormalTransistorPmos: -3.50179e+07 muA
** DiodeTransistorPmos: -3.45859e+07 muA
** NormalTransistorNmos: 3.45851e+07 muA
** NormalTransistorNmos: 3.45861e+07 muA
** DiodeTransistorNmos: 1.85841e+07 muA
** DiodeTransistorNmos: 5.44991e+07 muA
** DiodeTransistorPmos: -1.00311e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.23101  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.915001  V
** inSourceTransconductanceComplementarySecondStage: 0.637001  V
** innerComplementarySecondStage: 4.18901  V
** inputVoltageBiasXXnXX0: 0.555001  V
** out: 2.5  V
** outFirstStage: 0.637001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40001  V
** sourceTransconductance: 3.24401  V
** innerStageBias: 4.65301  V
** innerTransconductance: 0.232001  V
** inner: 0.232001  V


.END