** Name: two_stage_single_output_op_amp_74_1

.MACRO two_stage_single_output_op_amp_74_1 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=78e-6
mMainBias2 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=10e-6 W=19e-6
mFoldedCascodeFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=67e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=63e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=82e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=78e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=24e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=24e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=67e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=19e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=301e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=8e-6 W=57e-6
mMainBias13 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=302e-6
mMainBias14 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=370e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=193e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=584e-6
mFoldedCascodeFirstStageLoad19 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=193e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.30001e-12
.EOM two_stage_single_output_op_amp_74_1

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 9.13601 mW
** Area: 14272 (mu_m)^2
** Transit frequency: 4.56301 MHz
** Transit frequency with error factor: 4.5632 MHz
** Slew rate: 5.54836 V/mu_s
** Phase margin: 60.1606°
** CMRR: 139 dB
** VoutMax: 4.64001 V
** VoutMin: 0.570001 V
** VcmMax: 5.04001 V
** VcmMin: 1.53001 V


** Expected Currents: 
** NormalTransistorNmos: 1.59916e+08 muA
** NormalTransistorNmos: 1.92269e+08 muA
** NormalTransistorPmos: -2.97139e+07 muA
** NormalTransistorPmos: -4.71229e+07 muA
** NormalTransistorPmos: -2.97129e+07 muA
** NormalTransistorPmos: -4.71219e+07 muA
** NormalTransistorNmos: 2.97131e+07 muA
** NormalTransistorNmos: 2.97121e+07 muA
** DiodeTransistorNmos: 2.97131e+07 muA
** NormalTransistorNmos: 3.48161e+07 muA
** DiodeTransistorNmos: 3.48171e+07 muA
** NormalTransistorNmos: 1.74081e+07 muA
** NormalTransistorNmos: 1.74081e+07 muA
** NormalTransistorNmos: 1.37087e+09 muA
** NormalTransistorPmos: -1.37086e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.59915e+08 muA
** DiodeTransistorPmos: -1.92268e+08 muA


** Expected Voltages: 
** ibias: 1.30601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.976001  V
** outSourceVoltageBiasXXnXX1: 0.654001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.07201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** out1: 1.18101  V
** sourceGCC1: 4.43501  V
** sourceGCC2: 4.43501  V
** sourceTransconductance: 1.86801  V
** inner: 0.651001  V


.END