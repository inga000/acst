** Name: two_stage_single_output_op_amp_4_2

.MACRO two_stage_single_output_op_amp_4_2 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=3e-6 W=19e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=30e-6
mSecondStage1StageBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=21e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=15e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=3e-6 W=30e-6
mSecondStage1Transconductor6 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=133e-6
mSecondStage1Transconductor7 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=301e-6
mSimpleFirstStageLoad8 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=3e-6 W=19e-6
mSimpleFirstStageTransconductor9 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=7e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=96e-6
mMainBias11 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=288e-6
mSecondStage1StageBias12 out ibias sourcePmos sourcePmos pmos4 L=6e-6 W=535e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=7e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_4_2

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 3.21901 mW
** Area: 8467 (mu_m)^2
** Transit frequency: 3.18601 MHz
** Transit frequency with error factor: 3.17569 MHz
** Slew rate: 14.4502 V/mu_s
** Phase margin: 63.0254°
** CMRR: 89 dB
** negPSRR: 89 dB
** posPSRR: 110 dB
** VoutMax: 4.53001 V
** VoutMin: 0.740001 V
** VcmMax: 3.24001 V
** VcmMin: 0.690001 V


** Expected Currents: 
** NormalTransistorPmos: -1.95485e+08 muA
** DiodeTransistorNmos: 3.25801e+07 muA
** DiodeTransistorNmos: 3.25791e+07 muA
** NormalTransistorNmos: 3.25801e+07 muA
** NormalTransistorNmos: 3.25791e+07 muA
** NormalTransistorPmos: -6.51619e+07 muA
** NormalTransistorPmos: -3.25809e+07 muA
** NormalTransistorPmos: -3.25809e+07 muA
** NormalTransistorNmos: 3.63144e+08 muA
** NormalTransistorNmos: 3.63143e+08 muA
** NormalTransistorPmos: -3.63143e+08 muA
** DiodeTransistorNmos: 1.95486e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 3.96101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.14401  V
** out: 2.5  V
** outFirstStage: 0.878001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 1.25201  V
** innerSourceLoad1: 0.601001  V
** innerTransistorStack2Load1: 0.600001  V
** sourceTransconductance: 3.78301  V
** innerTransconductance: 0.473001  V


.END