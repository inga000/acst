** Name: two_stage_single_output_op_amp_110_1

.MACRO two_stage_single_output_op_amp_110_1 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=224e-6
m2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=96e-6
m3 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=8e-6 W=96e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=12e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=163e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=225e-6
m7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=5e-6
m8 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=327e-6
m9 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=8e-6 W=96e-6
m10 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=269e-6
m11 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=203e-6
m12 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=96e-6
m13 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=370e-6
m14 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=6e-6
m15 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=73e-6
m16 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=225e-6
m17 FirstStageYinnerOutputLoad2 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=6e-6
m18 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=55e-6
m19 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=6e-6 W=55e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=163e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_110_1

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 2.84301 mW
** Area: 13395 (mu_m)^2
** Transit frequency: 4.28401 MHz
** Transit frequency with error factor: 4.28432 MHz
** Slew rate: 12.7041 V/mu_s
** Phase margin: 63.0254°
** CMRR: 131 dB
** VoutMax: 4.63001 V
** VoutMin: 0.300001 V
** VcmMax: 3.18001 V
** VcmMin: 1.20001 V


** Expected Currents: 
** NormalTransistorNmos: 7.31931e+07 muA
** NormalTransistorNmos: 5.52981e+07 muA
** NormalTransistorPmos: -6.13109e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** DiodeTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** DiodeTransistorNmos: 2.28561e+07 muA
** NormalTransistorPmos: -1.01015e+08 muA
** DiodeTransistorPmos: -1.01016e+08 muA
** NormalTransistorPmos: -2.28579e+07 muA
** NormalTransistorPmos: -2.28579e+07 muA
** NormalTransistorNmos: 3.13063e+08 muA
** NormalTransistorPmos: -3.13062e+08 muA
** DiodeTransistorNmos: 6.13101e+07 muA
** DiodeTransistorPmos: -7.31939e+07 muA
** NormalTransistorPmos: -7.31949e+07 muA
** DiodeTransistorPmos: -5.52989e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.06101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outInputVoltageBiasXXpXX1: 3.55401  V
** outSourceVoltageBiasXXpXX1: 4.27701  V
** outVoltageBiasXXnXX0: 0.555001  V
** outVoltageBiasXXpXX2: 1.76501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.43601  V
** innerOutputLoad2: 1.11001  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.555001  V
** sourceGCC1: 2.98501  V
** sourceGCC2: 2.97901  V
** inner: 4.27601  V


.END