** Name: two_stage_single_output_op_amp_64_9

.MACRO two_stage_single_output_op_amp_64_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=147e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=40e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=333e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=122e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=6e-6 W=169e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=6e-6 W=93e-6
mMainBias7 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=57e-6
mFoldedCascodeFirstStageStageBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=125e-6
mFoldedCascodeFirstStageLoad9 FirstStageYinnerOutputLoad2 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=38e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=50e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=50e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=40e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=333e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=38e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=6e-6 W=93e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=58e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=58e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=125e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=57e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=403e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=253e-6
mFoldedCascodeFirstStageLoad22 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=169e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=433e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_64_9

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 4.32901 mW
** Area: 13494 (mu_m)^2
** Transit frequency: 2.83401 MHz
** Transit frequency with error factor: 2.83405 MHz
** Slew rate: 3.97006 V/mu_s
** Phase margin: 65.8902°
** CMRR: 140 dB
** VoutMax: 4.25 V
** VoutMin: 0.700001 V
** VcmMax: 3.15001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorPmos: -7.61869e+07 muA
** NormalTransistorPmos: -7.04409e+07 muA
** NormalTransistorNmos: 1.80941e+07 muA
** NormalTransistorNmos: 2.92141e+07 muA
** NormalTransistorNmos: 1.80941e+07 muA
** NormalTransistorNmos: 2.92141e+07 muA
** DiodeTransistorPmos: -1.80949e+07 muA
** DiodeTransistorPmos: -1.80959e+07 muA
** NormalTransistorPmos: -1.80949e+07 muA
** NormalTransistorPmos: -1.80959e+07 muA
** NormalTransistorPmos: -2.22409e+07 muA
** DiodeTransistorPmos: -2.22399e+07 muA
** NormalTransistorPmos: -1.11209e+07 muA
** NormalTransistorPmos: -1.11209e+07 muA
** NormalTransistorNmos: 6.40647e+08 muA
** DiodeTransistorNmos: 6.40646e+08 muA
** NormalTransistorPmos: -6.40646e+08 muA
** DiodeTransistorNmos: 7.61861e+07 muA
** NormalTransistorNmos: 7.61861e+07 muA
** DiodeTransistorNmos: 7.04401e+07 muA
** DiodeTransistorNmos: 7.04411e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.42601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.12601  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.571001  V
** outSourceVoltageBiasXXpXX1: 4.21401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 3.42601  V
** innerTransistorStack1Load2: 4.18001  V
** innerTransistorStack2Load2: 4.17901  V
** sourceGCC1: 0.571001  V
** sourceGCC2: 0.571001  V
** sourceTransconductance: 3.33701  V
** inner: 0.555001  V
** inner: 4.21101  V


.END