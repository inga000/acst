.suckt  symmetrical_op_amp200 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_MainBias_1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_2 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_3 out1FirstStage out1FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m_Symmetrical_FirstStage_Load_4 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Load_5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_Symmetrical_FirstStage_Load_6 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_StageBias_7 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_Symmetrical_FirstStage_StageBias_8 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Transconductor_9 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_Symmetrical_FirstStage_Transconductor_10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_StageBias_11 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m_Symmetrical_SecondStage1_StageBias_12 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_Transconductor_13 out out1FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m_Symmetrical_SecondStage1_Transconductor_14 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_15 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_16 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_17 innerComplementarySecondStage inSourceTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_MainBias_19 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_20 ibias ibias sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_21 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end symmetrical_op_amp200

