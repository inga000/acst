** Name: one_stage_single_output_op_amp67

.MACRO one_stage_single_output_op_amp67 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=53e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=176e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=6e-6 W=129e-6
mFoldedCascodeFirstStageLoad4 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=129e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=13e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerOutputLoad2 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=22e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=144e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=144e-6
mFoldedCascodeFirstStageLoad10 out inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=22e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=185e-6
mFoldedCascodeFirstStageLoad12 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=129e-6
mFoldedCascodeFirstStageTransconductor13 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=456e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=456e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=363e-6
mMainBias16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=333e-6
mFoldedCascodeFirstStageLoad17 out FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=129e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp67

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 4.51901 mW
** Area: 5353 (mu_m)^2
** Transit frequency: 9.75201 MHz
** Transit frequency with error factor: 9.75216 MHz
** Slew rate: 9.07423 V/mu_s
** Phase margin: 89.3815°
** CMRR: 127 dB
** VoutMax: 3.35001 V
** VoutMin: 0.870001 V
** VcmMax: 3.32001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -3.35214e+08 muA
** NormalTransistorNmos: 1.81799e+08 muA
** NormalTransistorNmos: 2.74268e+08 muA
** NormalTransistorNmos: 1.81799e+08 muA
** NormalTransistorNmos: 2.74268e+08 muA
** DiodeTransistorPmos: -1.81798e+08 muA
** NormalTransistorPmos: -1.81799e+08 muA
** NormalTransistorPmos: -1.81798e+08 muA
** DiodeTransistorPmos: -1.81799e+08 muA
** NormalTransistorPmos: -1.8494e+08 muA
** NormalTransistorPmos: -1.84941e+08 muA
** NormalTransistorPmos: -9.24699e+07 muA
** NormalTransistorPmos: -9.24699e+07 muA
** DiodeTransistorNmos: 3.35215e+08 muA
** DiodeTransistorNmos: 3.35216e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.42701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.23201  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 2.78201  V
** innerStageBias: 4.16001  V
** innerTransistorStack1Load2: 4.03101  V
** innerTransistorStack2Load2: 4.03701  V
** sourceGCC1: 0.513001  V
** sourceGCC2: 0.513001  V
** sourceTransconductance: 3.21401  V


.END