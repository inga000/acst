** Name: two_stage_single_output_op_amp_206_8

.MACRO two_stage_single_output_op_amp_206_8 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=54e-6
m2 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=8e-6 W=8e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=43e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
m5 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=12e-6
m6 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
m7 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=41e-6
m8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=9e-6
m9 out outInputVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=8e-6 W=69e-6
m10 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=1e-6 W=12e-6
m11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=19e-6
m12 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=19e-6
m13 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
m14 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=43e-6
m15 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=69e-6
m16 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=54e-6
m17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
m18 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=598e-6
m19 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=20e-6
m20 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=42e-6
m21 FirstStageYinnerOutputLoad1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=598e-6
m22 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=262e-6
m23 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=262e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_206_8

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 5.48901 mW
** Area: 10605 (mu_m)^2
** Transit frequency: 2.56501 MHz
** Transit frequency with error factor: 2.56104 MHz
** Slew rate: 3.78896 V/mu_s
** Phase margin: 61.3065°
** CMRR: 122 dB
** VoutMax: 4.25 V
** VoutMin: 1.90001 V
** VcmMax: 4.57001 V
** VcmMin: 1.44001 V


** Expected Currents: 
** NormalTransistorPmos: -2.23999e+07 muA
** NormalTransistorPmos: -4.71449e+07 muA
** DiodeTransistorNmos: 2.87868e+08 muA
** NormalTransistorNmos: 2.87869e+08 muA
** NormalTransistorNmos: 2.8787e+08 muA
** DiodeTransistorNmos: 2.87869e+08 muA
** NormalTransistorPmos: -2.9676e+08 muA
** NormalTransistorPmos: -2.96759e+08 muA
** NormalTransistorPmos: -2.9676e+08 muA
** NormalTransistorPmos: -2.96759e+08 muA
** NormalTransistorNmos: 1.77851e+07 muA
** DiodeTransistorNmos: 1.77841e+07 muA
** NormalTransistorNmos: 8.89301e+06 muA
** NormalTransistorNmos: 8.89301e+06 muA
** NormalTransistorNmos: 4.14834e+08 muA
** NormalTransistorNmos: 4.14833e+08 muA
** NormalTransistorPmos: -4.14833e+08 muA
** DiodeTransistorNmos: 2.23991e+07 muA
** NormalTransistorNmos: 2.23981e+07 muA
** DiodeTransistorNmos: 4.71441e+07 muA
** DiodeTransistorNmos: 4.71451e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.20401  V
** outInputVoltageBiasXXnXX2: 2.30301  V
** outSourceVoltageBiasXXnXX1: 0.602001  V
** outSourceVoltageBiasXXnXX2: 1.15501  V
** outSourceVoltageBiasXXpXX1: 3.93501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.09501  V
** innerSourceLoad1: 1.15501  V
** innerTransistorStack1Load1: 1.15601  V
** innerTransistorStack1Load2: 4.03301  V
** innerTransistorStack2Load2: 4.03301  V
** sourceTransconductance: 1.85901  V
** innerStageBias: 1.14801  V
** inner: 0.601001  V


.END