.suckt  complementary_op_amp15 ibias in1 in2 out sourceNmos sourcePmos
m_Complementary_MainBias_1 inputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_MainBias_2 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_Complementary_MainBias_3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_4 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m_Complementary_FirstStage_Load_5 FirstStageYinnerTransistorStack1LoadPmos FirstStageYout1 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_6 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m_Complementary_FirstStage_Load_7 FirstStageYinnerTransistorStack2LoadPmos FirstStageYout1 sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m_Complementary_FirstStage_Load_9 FirstStageYinnerTransistorStack1LoadNmos FirstStageYout1 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_10 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m_Complementary_FirstStage_Load_11 FirstStageYinnerTransistorStack2LoadNmos FirstStageYout1 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_12 FirstStageYsourceTransconductanceNmos outVoltageBiasXXnXX1 FirstStageYinnerStageBiasNmos FirstStageYinnerStageBiasNmos nmos
m_Complementary_FirstStage_StageBias_13 FirstStageYinnerStageBiasNmos inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_14 FirstStageYsourceTransconductancePmos inputVoltageBiasXXpXX1 FirstStageYinnerStageBiasPmos FirstStageYinnerStageBiasPmos pmos
m_Complementary_FirstStage_StageBias_15 FirstStageYinnerStageBiasPmos ibias sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Transconductor_16 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_17 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_18 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m_Complementary_FirstStage_Transconductor_19 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c_Complementary_Load_Capacitor_1 out sourceNmos 
m_Complementary_MainBias_20 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_MainBias_21 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_MainBias_22 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_Complementary_MainBias_23 ibias ibias sourcePmos sourcePmos pmos
.end complementary_op_amp15

