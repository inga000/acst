** Name: two_stage_single_output_op_amp_6_4

.MACRO two_stage_single_output_op_amp_6_4 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=15e-6
m2 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=279e-6
m3 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=1e-6 W=13e-6
m4 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=23e-6
m6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=16e-6
m7 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=104e-6
m8 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=1e-6 W=13e-6
m9 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=408e-6
m10 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
m11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=170e-6
m12 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=267e-6
m13 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=254e-6
m14 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=600e-6
m15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=15e-6
m16 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=15e-6
m17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=134e-6
m18 SecondStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=600e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_6_4

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 3.65401 mW
** Area: 9821 (mu_m)^2
** Transit frequency: 2.81301 MHz
** Transit frequency with error factor: 2.80427 MHz
** Slew rate: 10.5423 V/mu_s
** Phase margin: 64.7443°
** CMRR: 92 dB
** negPSRR: 85 dB
** posPSRR: 88 dB
** VoutMax: 4.57001 V
** VoutMin: 0.75 V
** VcmMax: 3.43001 V
** VcmMin: 0.570001 V


** Expected Currents: 
** NormalTransistorNmos: 1.62454e+08 muA
** NormalTransistorPmos: -1.12237e+08 muA
** NormalTransistorPmos: -1.1692e+08 muA
** DiodeTransistorNmos: 2.96051e+07 muA
** NormalTransistorNmos: 2.96041e+07 muA
** NormalTransistorNmos: 2.96051e+07 muA
** DiodeTransistorNmos: 2.96041e+07 muA
** NormalTransistorPmos: -5.92119e+07 muA
** NormalTransistorPmos: -2.96059e+07 muA
** NormalTransistorPmos: -2.96059e+07 muA
** NormalTransistorNmos: 2.59879e+08 muA
** NormalTransistorNmos: 2.59878e+08 muA
** NormalTransistorPmos: -2.59878e+08 muA
** NormalTransistorPmos: -2.59879e+08 muA
** DiodeTransistorNmos: 1.12238e+08 muA
** DiodeTransistorNmos: 1.16921e+08 muA
** DiodeTransistorPmos: -1.62453e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.16501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.559001  V
** inputVoltageBiasXXnXX1: 1.15201  V
** out: 2.5  V
** outFirstStage: 0.733001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 1.13801  V
** innerTransistorStack1Load1: 0.569001  V
** innerTransistorStack2Load1: 0.569001  V
** sourceTransconductance: 3.80401  V
** innerStageBias: 4.40501  V
** innerTransconductance: 0.328001  V


.END