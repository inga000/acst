** Name: two_stage_single_output_op_amp_74_10

.MACRO two_stage_single_output_op_amp_74_10 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=129e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=19e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=498e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=129e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=27e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=8e-6 W=27e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=498e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=19e-6
mSecondStage1StageBias12 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=600e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=7e-6 W=480e-6
mMainBias14 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=18e-6
mMainBias15 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=519e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=476e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=476e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=389e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=600e-6
mFoldedCascodeFirstStageLoad21 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=519e-6
mMainBias22 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 13.1001e-12
.EOM two_stage_single_output_op_amp_74_10

** Expected Performance Values: 
** Gain: 117 dB
** Power consumption: 9.41201 mW
** Area: 14993 (mu_m)^2
** Transit frequency: 5.11301 MHz
** Transit frequency with error factor: 5.11304 MHz
** Slew rate: 24.1137 V/mu_s
** Phase margin: 60.1606°
** CMRR: 126 dB
** VoutMax: 4.25 V
** VoutMin: 0.220001 V
** VcmMax: 5.17001 V
** VcmMin: 1.91001 V


** Expected Currents: 
** NormalTransistorNmos: 2.53821e+07 muA
** NormalTransistorNmos: 1.13401e+07 muA
** NormalTransistorPmos: -1.22979e+07 muA
** NormalTransistorPmos: -3.21886e+08 muA
** NormalTransistorPmos: -4.82828e+08 muA
** NormalTransistorPmos: -3.21889e+08 muA
** NormalTransistorPmos: -4.82833e+08 muA
** NormalTransistorNmos: 3.21889e+08 muA
** NormalTransistorNmos: 3.2189e+08 muA
** DiodeTransistorNmos: 3.21889e+08 muA
** NormalTransistorNmos: 3.21886e+08 muA
** DiodeTransistorNmos: 3.21885e+08 muA
** NormalTransistorNmos: 1.60944e+08 muA
** NormalTransistorNmos: 1.60944e+08 muA
** NormalTransistorNmos: 8.57684e+08 muA
** NormalTransistorPmos: -8.57683e+08 muA
** NormalTransistorPmos: -8.57684e+08 muA
** DiodeTransistorNmos: 1.22971e+07 muA
** NormalTransistorNmos: 1.22961e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.53829e+07 muA
** DiodeTransistorPmos: -1.13409e+07 muA


** Expected Voltages: 
** ibias: 0.629001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.08401  V
** outInputVoltageBiasXXnXX1: 1.15801  V
** outSourceVoltageBiasXXnXX1: 0.579001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.19701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.647001  V
** out1: 1.28701  V
** sourceGCC1: 4.51301  V
** sourceGCC2: 4.51301  V
** sourceTransconductance: 1.34501  V
** innerTransconductance: 4.64801  V
** inner: 0.578001  V


.END