** Name: two_stage_single_output_op_amp_45_2

.MACRO two_stage_single_output_op_amp_45_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=13e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=17e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=10e-6 W=34e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
m6 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=66e-6
m7 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=31e-6
m8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=25e-6
m9 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=25e-6
m10 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=145e-6
m11 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=145e-6
m12 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=180e-6
m13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=10e-6 W=521e-6
m14 out ibias sourcePmos sourcePmos pmos4 L=10e-6 W=479e-6
m15 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=36e-6
m16 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=10e-6 W=22e-6
m17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=53e-6
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=8e-6
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=8e-6
m20 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=10e-6 W=153e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_45_2

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 2.29401 mW
** Area: 14903 (mu_m)^2
** Transit frequency: 2.85001 MHz
** Transit frequency with error factor: 2.84944 MHz
** Slew rate: 5.8222 V/mu_s
** Phase margin: 65.3172°
** CMRR: 132 dB
** VoutMax: 4.59001 V
** VoutMin: 0.5 V
** VcmMax: 3.47001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.53821e+07 muA
** NormalTransistorPmos: -1.53187e+08 muA
** NormalTransistorPmos: -6.47699e+06 muA
** NormalTransistorNmos: 3.23601e+07 muA
** NormalTransistorNmos: 5.52351e+07 muA
** NormalTransistorNmos: 3.23601e+07 muA
** NormalTransistorNmos: 5.52351e+07 muA
** DiodeTransistorPmos: -3.23609e+07 muA
** NormalTransistorPmos: -3.23609e+07 muA
** NormalTransistorPmos: -3.23609e+07 muA
** NormalTransistorPmos: -4.57469e+07 muA
** NormalTransistorPmos: -2.28739e+07 muA
** NormalTransistorPmos: -2.28739e+07 muA
** NormalTransistorNmos: 1.43223e+08 muA
** NormalTransistorNmos: 1.43222e+08 muA
** NormalTransistorPmos: -1.43222e+08 muA
** DiodeTransistorNmos: 1.53188e+08 muA
** DiodeTransistorNmos: 6.47601e+06 muA
** DiodeTransistorPmos: -2.53829e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.02901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.930001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.573001  V
** outVoltageBiasXXnXX2: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.56601  V
** out1: 4.25101  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.62701  V
** innerTransconductance: 0.193001  V


.END