** Name: two_stage_single_output_op_amp_71_7

.MACRO two_stage_single_output_op_amp_71_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=22e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=67e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=221e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=21e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=21e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=8e-6 W=46e-6
mSecondStage1StageBias10 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=265e-6
mFoldedCascodeFirstStageLoad11 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=22e-6
mFoldedCascodeFirstStageLoad12 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=42e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mMainBias15 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=356e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=10e-6 W=600e-6
mFoldedCascodeFirstStageLoad17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=42e-6
mMainBias18 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=506e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_71_7

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 7.75001 mW
** Area: 9295 (mu_m)^2
** Transit frequency: 3.70001 MHz
** Transit frequency with error factor: 3.69451 MHz
** Slew rate: 3.77639 V/mu_s
** Phase margin: 60.7336°
** CMRR: 107 dB
** VoutMax: 4.25 V
** VoutMin: 0.230001 V
** VcmMax: 5.17001 V
** VcmMin: 1.42001 V


** Expected Currents: 
** NormalTransistorPmos: -3.60939e+08 muA
** NormalTransistorPmos: -5.07107e+08 muA
** NormalTransistorPmos: -1.70569e+07 muA
** NormalTransistorPmos: -2.63599e+07 muA
** NormalTransistorPmos: -1.70569e+07 muA
** NormalTransistorPmos: -2.63599e+07 muA
** DiodeTransistorNmos: 1.70561e+07 muA
** NormalTransistorNmos: 1.70561e+07 muA
** NormalTransistorNmos: 1.86031e+07 muA
** NormalTransistorNmos: 1.86021e+07 muA
** NormalTransistorNmos: 9.30201e+06 muA
** NormalTransistorNmos: 9.30201e+06 muA
** NormalTransistorNmos: 6.09204e+08 muA
** NormalTransistorPmos: -6.09203e+08 muA
** DiodeTransistorNmos: 3.6094e+08 muA
** DiodeTransistorNmos: 5.07108e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.11501  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.639001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.514001  V
** out1: 0.570001  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.91701  V


.END