.suckt  one_stage_fully_differential_op_amp8 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
m_FullyDifferential_MainBias_1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_3 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_Load_5 outFeedback outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_6 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_8 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX1 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackStage_Transconductor_10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FeedbackStage_Transconductor_13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FirstStage_Load_14 out1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m_FullyDifferential_FirstStage_Load_15 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_16 out2 outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m_FullyDifferential_FirstStage_Load_17 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_18 out1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m_FullyDifferential_FirstStage_Load_19 FirstStageYinnerTransistorStack1Load2 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_20 out2 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m_FullyDifferential_FirstStage_Load_21 FirstStageYinnerTransistorStack2Load2 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_StageBias_22 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Transconductor_23 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_FullyDifferential_FirstStage_Transconductor_24 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_FullyDifferential_Load_Capacitor_1 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_2 out2 sourceNmos 
m_FullyDifferential_MainBias_25 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_26 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_27 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_28 ibias ibias sourcePmos sourcePmos pmos
.end one_stage_fully_differential_op_amp8

