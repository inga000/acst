** Name: two_stage_single_output_op_amp_138_3

.MACRO two_stage_single_output_op_amp_138_3 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=10e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
m3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=44e-6
m5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=86e-6
m6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=4e-6 W=86e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=192e-6
m8 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=61e-6
m9 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=135e-6
m10 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=113e-6
m11 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=392e-6
m12 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=392e-6
m13 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=3e-6 W=135e-6
m14 out outVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=6e-6 W=378e-6
m15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=86e-6
m16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=15e-6
m17 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=4e-6 W=86e-6
m18 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=15e-6
m19 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=91e-6
m20 SecondStageYinnerStageBias inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=372e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_138_3

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 4.74501 mW
** Area: 9449 (mu_m)^2
** Transit frequency: 3.43801 MHz
** Transit frequency with error factor: 3.42617 MHz
** Slew rate: 12.6173 V/mu_s
** Phase margin: 60.1606°
** CMRR: 93 dB
** VoutMax: 4.26001 V
** VoutMin: 0.340001 V
** VcmMax: 3.47001 V
** VcmMin: -0.149999 V


** Expected Currents: 
** NormalTransistorNmos: 7.44571e+07 muA
** NormalTransistorNmos: 3.99481e+07 muA
** DiodeTransistorPmos: -2.18297e+08 muA
** NormalTransistorPmos: -2.18297e+08 muA
** NormalTransistorPmos: -2.18297e+08 muA
** DiodeTransistorPmos: -2.18297e+08 muA
** NormalTransistorNmos: 2.56373e+08 muA
** NormalTransistorNmos: 2.56372e+08 muA
** NormalTransistorNmos: 2.56373e+08 muA
** NormalTransistorNmos: 2.56372e+08 muA
** NormalTransistorPmos: -7.61509e+07 muA
** NormalTransistorPmos: -3.80749e+07 muA
** NormalTransistorPmos: -3.80749e+07 muA
** NormalTransistorNmos: 3.11865e+08 muA
** NormalTransistorPmos: -3.11864e+08 muA
** NormalTransistorPmos: -3.11865e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.44579e+07 muA
** DiodeTransistorPmos: -3.99489e+07 muA


** Expected Voltages: 
** ibias: 1.15101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.21901  V
** out: 2.5  V
** outFirstStage: 0.746001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 3.68601  V
** innerTransistorStack1Load2: 0.486001  V
** innerTransistorStack2Load1: 3.68601  V
** innerTransistorStack2Load2: 0.486001  V
** out1: 2.37201  V
** sourceTransconductance: 3.81401  V
** innerStageBias: 4.77401  V


.END