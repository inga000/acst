** Name: two_stage_single_output_op_amp_24_5

.MACRO two_stage_single_output_op_amp_24_5 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=6e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=37e-6
m3 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=2e-6 W=12e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=69e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=403e-6
m6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=532e-6
m8 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=157e-6
m9 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=10e-6 W=130e-6
m10 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=157e-6
m11 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=156e-6
m12 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=156e-6
m13 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=2e-6 W=600e-6
m14 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=27e-6
m15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=299e-6
m16 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=17e-6
m17 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=299e-6
m18 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=403e-6
m19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=69e-6
m20 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=12e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.10001e-12
.EOM two_stage_single_output_op_amp_24_5

** Expected Performance Values: 
** Gain: 99 dB
** Power consumption: 4.57101 mW
** Area: 11664 (mu_m)^2
** Transit frequency: 11.6701 MHz
** Transit frequency with error factor: 11.6458 MHz
** Slew rate: 17.2763 V/mu_s
** Phase margin: 60.1606°
** CMRR: 97 dB
** negPSRR: 99 dB
** posPSRR: 171 dB
** VoutMax: 3.82001 V
** VoutMin: 0.150001 V
** VcmMax: 3.02001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 5.08041e+07 muA
** NormalTransistorPmos: -1.43659e+07 muA
** NormalTransistorPmos: -2.28169e+07 muA
** NormalTransistorNmos: 1.49577e+08 muA
** NormalTransistorNmos: 1.49576e+08 muA
** NormalTransistorNmos: 1.49577e+08 muA
** NormalTransistorNmos: 1.49576e+08 muA
** NormalTransistorPmos: -2.99154e+08 muA
** DiodeTransistorPmos: -2.99155e+08 muA
** NormalTransistorPmos: -1.49576e+08 muA
** NormalTransistorPmos: -1.49576e+08 muA
** NormalTransistorNmos: 5.07055e+08 muA
** NormalTransistorPmos: -5.07053e+08 muA
** DiodeTransistorPmos: -5.07052e+08 muA
** DiodeTransistorNmos: 1.43651e+07 muA
** DiodeTransistorNmos: 2.28161e+07 muA
** DiodeTransistorPmos: -5.08049e+07 muA
** NormalTransistorPmos: -5.08059e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.25701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.46401  V
** outSourceVoltageBiasXXpXX1: 4.23201  V
** outSourceVoltageBiasXXpXX2: 4.13001  V
** outVoltageBiasXXnXX0: 0.619001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.50501  V
** inner: 4.23001  V
** inner: 4.125  V


.END