** Name: two_stage_single_output_op_amp_52_5

.MACRO two_stage_single_output_op_amp_52_5 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=181e-6
m2 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=13e-6
m3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=3e-6 W=19e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=14e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=592e-6
m7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
m8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=181e-6
m9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=101e-6
m10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=101e-6
m11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=9e-6 W=305e-6
m12 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=65e-6
m13 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=582e-6
m14 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=547e-6
m15 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=35e-6
m16 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=57e-6
m17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=124e-6
m18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=124e-6
m19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=14e-6
m20 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=18e-6
m21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=592e-6
m22 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=57e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 18.1001e-12
.EOM two_stage_single_output_op_amp_52_5

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 9.07701 mW
** Area: 14934 (mu_m)^2
** Transit frequency: 12.1771 MHz
** Transit frequency with error factor: 12.1768 MHz
** Slew rate: 9.45948 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 3.14001 V
** VoutMin: 0.150001 V
** VcmMax: 4.78001 V
** VcmMin: 0.850001 V


** Expected Currents: 
** NormalTransistorNmos: 2.64751e+07 muA
** NormalTransistorNmos: 4.98291e+07 muA
** NormalTransistorPmos: -4.27119e+07 muA
** NormalTransistorPmos: -1.73638e+08 muA
** NormalTransistorPmos: -2.8899e+08 muA
** NormalTransistorPmos: -1.73639e+08 muA
** NormalTransistorPmos: -2.88991e+08 muA
** DiodeTransistorNmos: 1.73639e+08 muA
** NormalTransistorNmos: 1.7364e+08 muA
** NormalTransistorNmos: 1.73639e+08 muA
** NormalTransistorNmos: 2.30704e+08 muA
** NormalTransistorNmos: 1.15352e+08 muA
** NormalTransistorNmos: 1.15352e+08 muA
** NormalTransistorNmos: 1.1085e+09 muA
** NormalTransistorPmos: -1.10849e+09 muA
** DiodeTransistorPmos: -1.10849e+09 muA
** DiodeTransistorNmos: 4.27111e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.64759e+07 muA
** NormalTransistorPmos: -2.64769e+07 muA
** DiodeTransistorPmos: -4.98299e+07 muA
** DiodeTransistorPmos: -4.98309e+07 muA


** Expected Voltages: 
** ibias: 0.690001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.905001  V
** inputVoltageBiasXXpXX2: 2.57801  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.57201  V
** outSourceVoltageBiasXXpXX1: 3.78601  V
** outSourceVoltageBiasXXpXX2: 3.80801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.350001  V
** out1: 0.555001  V
** sourceGCC1: 3.85401  V
** sourceGCC2: 3.85401  V
** sourceTransconductance: 1.93001  V
** inner: 3.78401  V


.END