** Name: symmetrical_op_amp94

.MACRO symmetrical_op_amp94 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias2 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=79e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias4 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=10e-6
mSymmetricalFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=37e-6
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=37e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=87e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=87e-6
mSymmetricalFirstStageLoad9 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=32e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor10 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=2e-6 W=67e-6
mSecondStage1Transconductor11 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=67e-6
mSymmetricalFirstStageLoad12 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=32e-6
mSymmetricalFirstStageStageBias13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=550e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mSymmetricalFirstStageTransconductor15 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=19e-6
mSecondStage1StageBias16 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=187e-6
mSymmetricalFirstStageTransconductor17 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=19e-6
mMainBias18 out2FirstStage ibias sourcePmos sourcePmos pmos4 L=6e-6 W=172e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp94

** Expected Performance Values: 
** Gain: 95 dB
** Power consumption: 1.39901 mW
** Area: 5967 (mu_m)^2
** Transit frequency: 4.09201 MHz
** Transit frequency with error factor: 4.09224 MHz
** Slew rate: 8.31937 V/mu_s
** Phase margin: 85.3708°
** CMRR: 148 dB
** negPSRR: 47 dB
** posPSRR: 70 dB
** VoutMax: 3.65001 V
** VoutMin: 0.320001 V
** VcmMax: 3.91001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.18489e+07 muA
** NormalTransistorNmos: 3.54491e+07 muA
** NormalTransistorNmos: 3.54481e+07 muA
** NormalTransistorNmos: 3.54491e+07 muA
** NormalTransistorNmos: 3.54481e+07 muA
** NormalTransistorPmos: -7.08989e+07 muA
** NormalTransistorPmos: -3.54499e+07 muA
** NormalTransistorPmos: -3.54499e+07 muA
** NormalTransistorNmos: 8.34661e+07 muA
** NormalTransistorNmos: 8.34651e+07 muA
** NormalTransistorPmos: -8.34669e+07 muA
** NormalTransistorPmos: -8.34679e+07 muA
** DiodeTransistorPmos: -8.36839e+07 muA
** DiodeTransistorPmos: -8.36849e+07 muA
** NormalTransistorNmos: 8.36831e+07 muA
** NormalTransistorNmos: 8.36821e+07 muA
** DiodeTransistorNmos: 2.18481e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.22901  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 3.80901  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 2.55801  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.726001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.159001  V
** innerTransistorStack2Load1: 0.159001  V
** sourceTransconductance: 3.38601  V
** innerStageBias: 3.28001  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END