.suckt  two_stage_fully_differential_op_amp_21_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m2 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m5 outFeedback outFeedback sourcePmos sourcePmos pmos
m6 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m7 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m8 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m9 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m10 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m12 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m13 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m14 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m15 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m16 sourceTransconductance inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m17 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m18 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m19 out1 outVoltageBiasXXnXX2 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m20 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m21 out1 ibias SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m22 SecondStage1YinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m23 out2 outVoltageBiasXXnXX2 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m24 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m25 out2 ibias SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m26 SecondStage2YinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m27 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
m28 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m29 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m30 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m31 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_21_4

