** Name: two_stage_single_output_op_amp_36_9

.MACRO two_stage_single_output_op_amp_36_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=2e-6 W=5e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=5e-6 W=286e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=23e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=271e-6
mSimpleFirstStageLoad5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=67e-6
mSimpleFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=6e-6 W=63e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=298e-6
mSimpleFirstStageTransconductor8 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=40e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=23e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=286e-6
mMainBias11 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias12 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=92e-6
mSecondStage1StageBias13 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=271e-6
mSimpleFirstStageTransconductor14 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=40e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=6e-6 W=67e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=290e-6
mSimpleFirstStageLoad17 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=6e-6 W=63e-6
mMainBias18 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=5e-6 W=338e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_36_9

** Expected Performance Values: 
** Gain: 95 dB
** Power consumption: 4.77201 mW
** Area: 10998 (mu_m)^2
** Transit frequency: 3.96701 MHz
** Transit frequency with error factor: 3.96397 MHz
** Slew rate: 3.73844 V/mu_s
** Phase margin: 60.7336°
** CMRR: 107 dB
** negPSRR: 101 dB
** posPSRR: 95 dB
** VoutMax: 4.36001 V
** VoutMin: 0.840001 V
** VcmMax: 3.86001 V
** VcmMin: 1.38001 V


** Expected Currents: 
** NormalTransistorNmos: 1.85212e+08 muA
** NormalTransistorPmos: -2.0741e+08 muA
** DiodeTransistorPmos: -8.46699e+06 muA
** DiodeTransistorPmos: -8.46799e+06 muA
** NormalTransistorPmos: -8.46699e+06 muA
** NormalTransistorPmos: -8.46799e+06 muA
** NormalTransistorNmos: 1.69311e+07 muA
** DiodeTransistorNmos: 1.69301e+07 muA
** NormalTransistorNmos: 8.46601e+06 muA
** NormalTransistorNmos: 8.46601e+06 muA
** NormalTransistorNmos: 5.34767e+08 muA
** DiodeTransistorNmos: 5.34768e+08 muA
** NormalTransistorPmos: -5.34766e+08 muA
** DiodeTransistorNmos: 2.07411e+08 muA
** NormalTransistorNmos: 2.07411e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.85211e+08 muA


** Expected Voltages: 
** ibias: 1.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.02001  V
** out: 2.5  V
** outFirstStage: 3.79101  V
** outInputVoltageBiasXXnXX1: 1.22601  V
** outSourceVoltageBiasXXnXX1: 0.613001  V
** outSourceVoltageBiasXXnXX2: 0.622001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.22901  V
** innerTransistorStack2Load1: 4.22801  V
** out1: 3.45201  V
** sourceTransconductance: 1.94501  V
** inner: 0.613001  V
** inner: 0.619001  V


.END