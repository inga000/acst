** Name: symmetrical_op_amp118

.MACRO symmetrical_op_amp118 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=12e-6
m2 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
m3 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m4 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=38e-6
m5 innerComplementarySecondStage inStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
m6 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage nmos4 L=1e-6 W=31e-6
m7 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=38e-6
m8 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=4e-6 W=120e-6
m9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=4e-6 W=201e-6
m10 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=205e-6
m11 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=184e-6
m12 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=184e-6
m13 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=205e-6
m14 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=51e-6
m15 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=51e-6
m16 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=46e-6
m17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=46e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp118

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 2.12601 mW
** Area: 3091 (mu_m)^2
** Transit frequency: 7.38001 MHz
** Transit frequency with error factor: 7.38006 MHz
** Slew rate: 7.45518 V/mu_s
** Phase margin: 83.6519°
** CMRR: 144 dB
** negPSRR: 114 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 1.14001 V
** VcmMax: 4.81001 V
** VcmMin: 0.760001 V


** Expected Currents: 
** NormalTransistorNmos: 1.00565e+08 muA
** NormalTransistorPmos: -8.25559e+07 muA
** NormalTransistorPmos: -8.25569e+07 muA
** NormalTransistorPmos: -8.25559e+07 muA
** NormalTransistorPmos: -8.25569e+07 muA
** NormalTransistorNmos: 1.65111e+08 muA
** NormalTransistorNmos: 8.25551e+07 muA
** NormalTransistorNmos: 8.25551e+07 muA
** NormalTransistorNmos: 7.47281e+07 muA
** DiodeTransistorNmos: 7.47271e+07 muA
** NormalTransistorPmos: -7.47289e+07 muA
** NormalTransistorPmos: -7.47289e+07 muA
** NormalTransistorNmos: 7.47281e+07 muA
** NormalTransistorPmos: -7.47289e+07 muA
** NormalTransistorPmos: -7.47289e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.00564e+08 muA


** Expected Voltages: 
** ibias: 0.603001  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** inStageBiasComplementarySecondStage: 0.969001  V
** innerComplementarySecondStage: 1.54201  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.93401  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END