** Name: two_stage_single_output_op_amp_113_9

.MACRO two_stage_single_output_op_amp_113_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=10e-6 W=29e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=115e-6
mMainBias4 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=30e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=26e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mTelescopicFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=459e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=33e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=33e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=33e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias13 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=115e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=33e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=128e-6
mMainBias17 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=48e-6
mSecondStage1Transconductor18 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=446e-6
mTelescopicFirstStageLoad19 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=26e-6
mMainBias20 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=114e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.1001e-12
.EOM two_stage_single_output_op_amp_113_9

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 2.03401 mW
** Area: 9526 (mu_m)^2
** Transit frequency: 2.75201 MHz
** Transit frequency with error factor: 2.75087 MHz
** Slew rate: 7.26397 V/mu_s
** Phase margin: 60.1606°
** CMRR: 94 dB
** VoutMax: 4.74001 V
** VoutMin: 0.880001 V
** VcmMax: 4.43001 V
** VcmMin: 1.40001 V


** Expected Currents: 
** NormalTransistorNmos: 9.94601e+06 muA
** NormalTransistorPmos: -2.35399e+07 muA
** NormalTransistorPmos: -5.65749e+07 muA
** NormalTransistorNmos: 1.57141e+07 muA
** NormalTransistorNmos: 1.57141e+07 muA
** DiodeTransistorPmos: -1.57149e+07 muA
** NormalTransistorPmos: -1.57149e+07 muA
** NormalTransistorNmos: 8.80011e+07 muA
** NormalTransistorNmos: 8.80001e+07 muA
** NormalTransistorNmos: 1.57141e+07 muA
** NormalTransistorNmos: 1.57141e+07 muA
** NormalTransistorNmos: 2.75384e+08 muA
** DiodeTransistorNmos: 2.75383e+08 muA
** NormalTransistorPmos: -2.75383e+08 muA
** DiodeTransistorNmos: 2.35391e+07 muA
** NormalTransistorNmos: 2.35391e+07 muA
** DiodeTransistorNmos: 5.65741e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.94699e+06 muA


** Expected Voltages: 
** ibias: 1.16101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.28401  V
** inputVoltageBiasXXpXX0: 4.27001  V
** out: 2.5  V
** outFirstStage: 4.17201  V
** outSourceVoltageBiasXXnXX1: 0.642001  V
** outSourceVoltageBiasXXnXX3: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.470001  V
** out1: 4.17501  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.642001  V


.END