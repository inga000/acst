** Name: two_stage_single_output_op_amp_64_8

.MACRO two_stage_single_output_op_amp_64_8 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=56e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=53e-6
m3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=5e-6 W=57e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=153e-6
m5 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=72e-6
m6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=29e-6
m7 out outInputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=543e-6
m8 outFirstStage outInputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
m9 FirstStageYinnerOutputLoad2 outInputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
m10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
m11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=16e-6
m12 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=532e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=216e-6
m14 outFirstStage FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=72e-6
m15 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=600e-6
m16 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack1Load2 sourcePmos sourcePmos pmos4 L=2e-6 W=29e-6
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=113e-6
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=113e-6
m19 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=153e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=57e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_64_8

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 6.34601 mW
** Area: 8076 (mu_m)^2
** Transit frequency: 5.83301 MHz
** Transit frequency with error factor: 5.83306 MHz
** Slew rate: 4.21252 V/mu_s
** Phase margin: 64.1713°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.710001 V
** VcmMax: 3.26001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.06719e+08 muA
** NormalTransistorNmos: 1.90551e+07 muA
** NormalTransistorNmos: 3.26671e+07 muA
** NormalTransistorNmos: 1.90511e+07 muA
** NormalTransistorNmos: 3.26611e+07 muA
** DiodeTransistorPmos: -1.90539e+07 muA
** DiodeTransistorPmos: -1.90529e+07 muA
** NormalTransistorPmos: -1.90519e+07 muA
** NormalTransistorPmos: -1.90529e+07 muA
** NormalTransistorPmos: -2.72219e+07 muA
** DiodeTransistorPmos: -2.72209e+07 muA
** NormalTransistorPmos: -1.36109e+07 muA
** NormalTransistorPmos: -1.36109e+07 muA
** NormalTransistorNmos: 1.07711e+09 muA
** NormalTransistorNmos: 1.07711e+09 muA
** NormalTransistorPmos: -1.0771e+09 muA
** DiodeTransistorNmos: 1.0672e+08 muA
** DiodeTransistorNmos: 1.06721e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.42601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.11501  V
** outSourceVoltageBiasXXnXX1: 0.560001  V
** outSourceVoltageBiasXXpXX1: 4.21401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad2: 3.42801  V
** innerTransistorStack1Load2: 4.16401  V
** innerTransistorStack2Load2: 4.16401  V
** sourceGCC1: 0.560001  V
** sourceGCC2: 0.560001  V
** sourceTransconductance: 3.22801  V
** innerStageBias: 0.557001  V
** inner: 4.21101  V


.END