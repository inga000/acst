** Name: two_stage_single_output_op_amp_50_3

.MACRO two_stage_single_output_op_amp_50_3 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=77e-6
mMainBias2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=36e-6
mMainBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=36e-6
mFoldedCascodeFirstStageTransconductor5 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=62e-6
mFoldedCascodeFirstStageTransconductor6 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=6e-6 W=62e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=123e-6
mMainBias8 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=296e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=457e-6
mFoldedCascodeFirstStageLoad10 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=77e-6
mFoldedCascodeFirstStageLoad11 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=366e-6
mFoldedCascodeFirstStageLoad12 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mFoldedCascodeFirstStageLoad13 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=22e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
mSecondStage1StageBias15 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=329e-6
mFoldedCascodeFirstStageLoad16 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=366e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9e-12
.EOM two_stage_single_output_op_amp_50_3

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 6.28701 mW
** Area: 3886 (mu_m)^2
** Transit frequency: 8.98201 MHz
** Transit frequency with error factor: 8.96434 MHz
** Slew rate: 14.9091 V/mu_s
** Phase margin: 60.1606°
** CMRR: 104 dB
** VoutMax: 3.42001 V
** VoutMin: 0.150001 V
** VcmMax: 4.66001 V
** VcmMin: 0.870001 V


** Expected Currents: 
** NormalTransistorNmos: 3.65522e+08 muA
** NormalTransistorPmos: -1.48014e+08 muA
** NormalTransistorPmos: -2.23373e+08 muA
** NormalTransistorPmos: -1.48014e+08 muA
** NormalTransistorPmos: -2.23373e+08 muA
** DiodeTransistorNmos: 1.48015e+08 muA
** NormalTransistorNmos: 1.48015e+08 muA
** NormalTransistorNmos: 1.50722e+08 muA
** NormalTransistorNmos: 7.53601e+07 muA
** NormalTransistorNmos: 7.53601e+07 muA
** NormalTransistorNmos: 4.35208e+08 muA
** NormalTransistorPmos: -4.35207e+08 muA
** NormalTransistorPmos: -4.35208e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.65521e+08 muA
** DiodeTransistorPmos: -3.65521e+08 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 2.37201  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceGCC1: 3.08601  V
** sourceGCC2: 3.08601  V
** sourceTransconductance: 1.80101  V
** innerStageBias: 3.20701  V


.END