.suckt  two_stage_fully_differential_op_amp_1_1 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m2 outFeedback outFeedback sourceNmos sourceNmos nmos
m3 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m4 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m5 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m6 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m7 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m8 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m9 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m10 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m11 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m12 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m13 out2FirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m14 out1 out1FirstStage sourceNmos sourceNmos nmos
m15 out1 ibias sourcePmos sourcePmos pmos
m16 out2 out2FirstStage sourceNmos sourceNmos nmos
m17 out2 ibias sourcePmos sourcePmos pmos
m18 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_1_1

