** Name: two_stage_single_output_op_amp_23_5

.MACRO two_stage_single_output_op_amp_23_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=24e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=6e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=530e-6
mMainBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad7 FirstStageYinnerSourceLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=344e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=159e-6
mSimpleFirstStageLoad9 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=1e-6 W=159e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
mSimpleFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=344e-6
mMainBias12 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
mSimpleFirstStageTransconductor13 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=205e-6
mSimpleFirstStageStageBias14 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
mSimpleFirstStageStageBias15 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=408e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mSecondStage1StageBias17 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=530e-6
mSimpleFirstStageTransconductor18 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=205e-6
mMainBias19 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=118e-6
mMainBias20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=26e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9e-12
.EOM two_stage_single_output_op_amp_23_5

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 14.9681 mW
** Area: 7523 (mu_m)^2
** Transit frequency: 36.6381 MHz
** Transit frequency with error factor: 36.5894 MHz
** Slew rate: 66.3329 V/mu_s
** Phase margin: 60.1606°
** CMRR: 101 dB
** negPSRR: 100 dB
** posPSRR: 134 dB
** VoutMax: 3.07001 V
** VoutMin: 0.210001 V
** VcmMax: 3.06001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.53341e+07 muA
** NormalTransistorPmos: -1.19636e+08 muA
** NormalTransistorPmos: -2.63599e+07 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04163e+08 muA
** NormalTransistorNmos: 3.04164e+08 muA
** NormalTransistorNmos: 3.04163e+08 muA
** NormalTransistorPmos: -6.08327e+08 muA
** NormalTransistorPmos: -6.08326e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorPmos: -3.04163e+08 muA
** NormalTransistorNmos: 2.19386e+09 muA
** NormalTransistorPmos: -2.19385e+09 muA
** DiodeTransistorPmos: -2.19385e+09 muA
** DiodeTransistorNmos: 1.19637e+08 muA
** DiodeTransistorNmos: 2.63591e+07 muA
** DiodeTransistorPmos: -2.53349e+07 muA
** NormalTransistorPmos: -2.53349e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.612001  V
** outInputVoltageBiasXXpXX1: 2.50401  V
** outSourceVoltageBiasXXpXX1: 3.75201  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.827001  V
** outVoltageBiasXXnXX1: 0.759001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerStageBias: 4.25  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.35101  V
** inner: 3.75201  V


.END