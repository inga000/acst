.suckt  two_stage_single_output_op_amp_170_6 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_3 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_4 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_6 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_SingleOutput_FirstStage_Load_7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_8 FirstStageYinnerOutputLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m_SingleOutput_FirstStage_Load_9 FirstStageYinnerTransistorStack1Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m_SingleOutput_FirstStage_Load_11 FirstStageYinnerTransistorStack2Load2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_StageBias_12 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_SingleOutput_FirstStage_StageBias_13 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Transconductor_14 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_SingleOutput_FirstStage_Transconductor_15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_Transconductor_16 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_SingleOutput_SecondStage1_Transconductor_17 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_18 out ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m_SingleOutput_SecondStage1_StageBias_19 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_20 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_21 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_22 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_SingleOutput_MainBias_23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_24 ibias ibias VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m_SingleOutput_MainBias_25 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_170_6

