** Name: one_stage_single_output_op_amp110

.MACRO one_stage_single_output_op_amp110 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=16e-6
m2 FirstStageYinnerOutputLoad2 FirstStageYinnerOutputLoad2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=47e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=47e-6
m4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=20e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=192e-6
m6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=5e-6
m7 out FirstStageYinnerOutputLoad2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=47e-6
m8 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=9e-6 W=13e-6
m9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=47e-6
m10 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m11 out outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=5e-6 W=270e-6
m12 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=192e-6
m13 FirstStageYinnerOutputLoad2 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=5e-6 W=270e-6
m14 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=48e-6
m15 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=48e-6
m16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp110

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 0.617001 mW
** Area: 3987 (mu_m)^2
** Transit frequency: 3.16901 MHz
** Transit frequency with error factor: 3.16874 MHz
** Slew rate: 4.86868 V/mu_s
** Phase margin: 75.0575°
** CMRR: 149 dB
** VoutMax: 3.65001 V
** VoutMin: 0.740001 V
** VcmMax: 3.30001 V
** VcmMin: 0.810001 V


** Expected Currents: 
** NormalTransistorNmos: 4.54701e+06 muA
** NormalTransistorPmos: -5.60399e+06 muA
** NormalTransistorPmos: -4.66349e+07 muA
** NormalTransistorPmos: -4.66349e+07 muA
** DiodeTransistorNmos: 4.66341e+07 muA
** NormalTransistorNmos: 4.66331e+07 muA
** NormalTransistorNmos: 4.66341e+07 muA
** DiodeTransistorNmos: 4.66331e+07 muA
** NormalTransistorPmos: -9.78159e+07 muA
** DiodeTransistorPmos: -9.78149e+07 muA
** NormalTransistorPmos: -4.66339e+07 muA
** NormalTransistorPmos: -4.66339e+07 muA
** DiodeTransistorNmos: 5.60301e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -4.54799e+06 muA


** Expected Voltages: 
** ibias: 3.53501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX0: 0.597001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.26801  V
** outVoltageBiasXXpXX2: 2.23001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.29601  V
** innerOutputLoad2: 1.15001  V
** innerSourceLoad2: 0.592001  V
** innerTransistorStack1Load2: 0.592001  V
** sourceGCC1: 3.01401  V
** sourceGCC2: 3.01401  V
** inner: 4.26601  V


.END