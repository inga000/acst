** Name: two_stage_single_output_op_amp_143_9

.MACRO two_stage_single_output_op_amp_143_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=11e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=283e-6
m3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=31e-6
m4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=13e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=5e-6 W=80e-6
m6 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=283e-6
m7 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=7e-6 W=7e-6
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=43e-6
m9 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=13e-6
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=43e-6
m11 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=54e-6
m12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
m13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=387e-6
m14 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=384e-6
m15 outFirstStage ibias sourcePmos sourcePmos pmos4 L=5e-6 W=495e-6
m16 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=189e-6
m17 FirstStageYout1 ibias sourcePmos sourcePmos pmos4 L=5e-6 W=495e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 8e-12
.EOM two_stage_single_output_op_amp_143_9

** Expected Performance Values: 
** Gain: 81 dB
** Power consumption: 7.45501 mW
** Area: 12786 (mu_m)^2
** Transit frequency: 5.34401 MHz
** Transit frequency with error factor: 5.33191 MHz
** Slew rate: 5.03679 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 1.32001 V
** VcmMax: 5.22001 V
** VcmMin: 0.770001 V


** Expected Currents: 
** NormalTransistorPmos: -4.88549e+07 muA
** NormalTransistorPmos: -2.38269e+07 muA
** NormalTransistorNmos: 4.12891e+07 muA
** NormalTransistorNmos: 4.12881e+07 muA
** DiodeTransistorNmos: 4.12891e+07 muA
** NormalTransistorPmos: -6.17639e+07 muA
** NormalTransistorPmos: -6.17639e+07 muA
** NormalTransistorNmos: 4.09491e+07 muA
** NormalTransistorNmos: 2.04751e+07 muA
** NormalTransistorNmos: 2.04751e+07 muA
** NormalTransistorNmos: 1.27471e+09 muA
** DiodeTransistorNmos: 1.27471e+09 muA
** NormalTransistorPmos: -1.2747e+09 muA
** DiodeTransistorNmos: 4.88541e+07 muA
** NormalTransistorNmos: 4.88531e+07 muA
** DiodeTransistorNmos: 2.38261e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.73001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.865001  V
** outVoltageBiasXXnXX2: 0.617001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.989001  V
** out1: 2.09501  V
** sourceTransconductance: 1.94501  V
** inner: 0.865001  V


.END