** Name: two_stage_single_output_op_amp_62_7

.MACRO two_stage_single_output_op_amp_62_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=118e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=199e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=40e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=223e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=7e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=89e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=166e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=166e-6
mSecondStage1StageBias10 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=600e-6
mFoldedCascodeFirstStageLoad11 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=89e-6
mMainBias12 outVoltageBiasXXpXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=17e-6
mFoldedCascodeFirstStageLoad13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=199e-6
mFoldedCascodeFirstStageTransconductor14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=55e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=55e-6
mFoldedCascodeFirstStageStageBias16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=223e-6
mMainBias17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=242e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=507e-6
mFoldedCascodeFirstStageLoad20 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=7e-6 W=384e-6
mMainBias21 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=115e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 14.2001e-12
.EOM two_stage_single_output_op_amp_62_7

** Expected Performance Values: 
** Gain: 132 dB
** Power consumption: 2.99201 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 3.70001 MHz
** Transit frequency with error factor: 3.69978 MHz
** Slew rate: 3.92848 V/mu_s
** Phase margin: 60.1606°
** CMRR: 144 dB
** VoutMax: 4.81001 V
** VoutMin: 0.190001 V
** VcmMax: 3.23001 V
** VcmMin: -0.369999 V


** Expected Currents: 
** NormalTransistorNmos: 8.83801e+06 muA
** NormalTransistorPmos: -2.85859e+07 muA
** NormalTransistorPmos: -6.01329e+07 muA
** NormalTransistorNmos: 5.63301e+07 muA
** NormalTransistorNmos: 8.45921e+07 muA
** NormalTransistorNmos: 5.63291e+07 muA
** NormalTransistorNmos: 8.45921e+07 muA
** DiodeTransistorPmos: -5.63309e+07 muA
** NormalTransistorPmos: -5.63299e+07 muA
** NormalTransistorPmos: -5.63309e+07 muA
** NormalTransistorPmos: -5.65239e+07 muA
** DiodeTransistorPmos: -5.65229e+07 muA
** NormalTransistorPmos: -2.82619e+07 muA
** NormalTransistorPmos: -2.82619e+07 muA
** NormalTransistorNmos: 3.11598e+08 muA
** NormalTransistorPmos: -3.11597e+08 muA
** DiodeTransistorNmos: 2.85851e+07 muA
** DiodeTransistorNmos: 6.01321e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -8.83899e+06 muA


** Expected Voltages: 
** ibias: 3.39601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.596001  V
** out: 2.5  V
** outFirstStage: 4.25  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.989001  V
** outVoltageBiasXXpXX2: 3.73001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.53301  V
** out1: 4.25801  V
** sourceGCC1: 0.391001  V
** sourceGCC2: 0.391001  V
** sourceTransconductance: 3.23301  V
** inner: 4.19601  V


.END