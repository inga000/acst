** Name: symmetrical_op_amp55

.MACRO symmetrical_op_amp55 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=41e-6
mSecondStage1StageBias5 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=8e-6 W=43e-6
mSymmetricalFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=144e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=31e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=31e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=2e-6 W=11e-6
mSecondStage1Transconductor10 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=11e-6
mSymmetricalFirstStageStageBias11 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=144e-6
mMainBias12 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=41e-6
mMainBias13 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=314e-6
mSymmetricalFirstStageTransconductor14 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=82e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias15 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=8e-6 W=43e-6
mSecondStage1StageBias16 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=1e-6 W=81e-6
mSymmetricalFirstStageTransconductor17 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=82e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp55

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 1.15901 mW
** Area: 4223 (mu_m)^2
** Transit frequency: 5.11501 MHz
** Transit frequency with error factor: 5.11519 MHz
** Slew rate: 4.94252 V/mu_s
** Phase margin: 79.0682°
** CMRR: 145 dB
** negPSRR: 53 dB
** posPSRR: 68 dB
** VoutMax: 3.53001 V
** VoutMin: 0.600001 V
** VcmMax: 3.25 V
** VcmMin: 0.120001 V


** Expected Currents: 
** NormalTransistorPmos: -7.72119e+07 muA
** DiodeTransistorNmos: 1.77901e+07 muA
** DiodeTransistorNmos: 1.77901e+07 muA
** NormalTransistorPmos: -3.55819e+07 muA
** DiodeTransistorPmos: -3.55809e+07 muA
** NormalTransistorPmos: -1.77909e+07 muA
** NormalTransistorPmos: -1.77909e+07 muA
** NormalTransistorNmos: 4.94791e+07 muA
** NormalTransistorNmos: 4.94801e+07 muA
** NormalTransistorPmos: -4.94799e+07 muA
** DiodeTransistorPmos: -4.94809e+07 muA
** NormalTransistorPmos: -4.94819e+07 muA
** NormalTransistorNmos: 4.94811e+07 muA
** NormalTransistorNmos: 4.94801e+07 muA
** DiodeTransistorNmos: 7.72111e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40201  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 1.00601  V
** inSourceTransconductanceComplementarySecondStage: 0.681001  V
** inStageBiasComplementarySecondStage: 3.71501  V
** innerComplementarySecondStage: 2.96601  V
** out: 2.5  V
** outFirstStage: 0.681001  V
** outSourceVoltageBiasXXpXX1: 4.20201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.22001  V
** innerTransconductance: 0.276001  V
** inner: 0.276001  V
** inner: 4.19901  V


.END