.suckt  two_stage_single_output_op_amp_10_10 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad3 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mSimpleFirstStageLoad4 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos
mSimpleFirstStageStageBias5 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSimpleFirstStageTransconductor7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1StageBias8 out ibias sourceNmos sourceNmos nmos
mSecondStage1Transconductor9 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
mMainBias11 ibias ibias sourceNmos sourceNmos nmos
mMainBias12 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_10_10

