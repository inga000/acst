.suckt  symmetrical_op_amp58 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m3 outFirstStage outFirstStage sourcePmos sourcePmos pmos
m4 inTransconductanceComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m5 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m6 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos
m7 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m8 inTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c1 out sourceNmos 
m9 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
m10 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
m11 out outFirstStage sourcePmos sourcePmos pmos
m12 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
m13 innerComplementarySecondStage inTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
m14 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m15 ibias ibias sourceNmos sourceNmos nmos
m16 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end symmetrical_op_amp58

