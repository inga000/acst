** Name: two_stage_single_output_op_amp_137_1

.MACRO two_stage_single_output_op_amp_137_1 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
m2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=62e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=3e-6 W=62e-6
m5 outFirstStage outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
m6 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=565e-6
m7 FirstStageYout1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=83e-6
m8 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=3e-6 W=62e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=3e-6 W=62e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=87e-6
m11 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
m12 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
m13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=124e-6
m14 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=87e-6
Capacitor1 outFirstStage out 15.9001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_137_1

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 4.47601 mW
** Area: 4263 (mu_m)^2
** Transit frequency: 4.77001 MHz
** Transit frequency with error factor: 4.75432 MHz
** Slew rate: 4.61043 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** VoutMax: 4.82001 V
** VoutMin: 0.150001 V
** VcmMax: 4.10001 V
** VcmMin: -0.149999 V


** Expected Currents: 
** NormalTransistorPmos: -2.33179e+07 muA
** DiodeTransistorPmos: -2.09836e+08 muA
** NormalTransistorPmos: -2.09836e+08 muA
** NormalTransistorPmos: -2.09836e+08 muA
** DiodeTransistorPmos: -2.09836e+08 muA
** NormalTransistorNmos: 2.46623e+08 muA
** NormalTransistorNmos: 2.46623e+08 muA
** NormalTransistorPmos: -7.35729e+07 muA
** NormalTransistorPmos: -3.67859e+07 muA
** NormalTransistorPmos: -3.67859e+07 muA
** NormalTransistorNmos: 3.58735e+08 muA
** NormalTransistorPmos: -3.58734e+08 muA
** DiodeTransistorNmos: 2.33191e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX1: 0.822001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.68601  V
** innerTransistorStack1Load1: 3.68601  V
** out1: 2.37201  V
** sourceTransconductance: 3.21801  V


.END