.suckt  complementary_op_amp23 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m3 FirstStageYout1 ibias FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m4 FirstStageYinnerTransistorStack1LoadNmos outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m5 out ibias FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m6 FirstStageYinnerTransistorStack2LoadNmos outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m7 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1LoadPmos FirstStageYinnerTransistorStack1LoadPmos pmos
m8 FirstStageYinnerTransistorStack1LoadPmos FirstStageYout1 sourcePmos sourcePmos pmos
m9 out outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m10 FirstStageYinnerTransistorStack2LoadPmos FirstStageYout1 sourcePmos sourcePmos pmos
m11 FirstStageYsourceTransconductanceNmos ibias FirstStageYinnerStageBiasNmos FirstStageYinnerStageBiasNmos nmos
m12 FirstStageYinnerStageBiasNmos outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m13 FirstStageYsourceTransconductancePmos outVoltageBiasXXpXX1 FirstStageYinnerStageBiasPmos FirstStageYinnerStageBiasPmos pmos
m14 FirstStageYinnerStageBiasPmos outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m15 FirstStageYinnerTransistorStack1LoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m16 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m17 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m18 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c1 out sourceNmos 
m19 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m20 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m21 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m22 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end complementary_op_amp23

