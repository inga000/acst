** Name: one_stage_single_output_op_amp122

.MACRO one_stage_single_output_op_amp122 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=5e-6
mTelescopicFirstStageStageBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=95e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=20e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=325e-6
mTelescopicFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=107e-6
mTelescopicFirstStageTransconductor7 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=215e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=215e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
mTelescopicFirstStageLoad11 out outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=107e-6
mMainBias12 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=35e-6
mTelescopicFirstStageStageBias13 sourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=95e-6
mTelescopicFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
mTelescopicFirstStageLoad15 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
mTelescopicFirstStageLoad16 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=84e-6
mTelescopicFirstStageLoad17 out inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=84e-6
mMainBias18 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=3e-6 W=244e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp122

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 1.41301 mW
** Area: 5915 (mu_m)^2
** Transit frequency: 7.22001 MHz
** Transit frequency with error factor: 7.22003 MHz
** Slew rate: 9.34541 V/mu_s
** Phase margin: 85.3708°
** CMRR: 144 dB
** VoutMax: 4.41001 V
** VoutMin: 1.14001 V
** VcmMax: 4.97001 V
** VcmMin: 1.39001 V


** Expected Currents: 
** NormalTransistorNmos: 6.90661e+07 muA
** NormalTransistorNmos: 1.61051e+07 muA
** NormalTransistorPmos: -5.09639e+07 muA
** NormalTransistorNmos: 6.82491e+07 muA
** NormalTransistorNmos: 6.82491e+07 muA
** NormalTransistorPmos: -6.825e+07 muA
** NormalTransistorPmos: -6.82509e+07 muA
** NormalTransistorPmos: -6.825e+07 muA
** NormalTransistorPmos: -6.82509e+07 muA
** NormalTransistorNmos: 1.87465e+08 muA
** DiodeTransistorNmos: 1.87466e+08 muA
** NormalTransistorNmos: 6.82501e+07 muA
** NormalTransistorNmos: 6.82501e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 5.09631e+07 muA
** DiodeTransistorPmos: -6.90669e+07 muA
** DiodeTransistorPmos: -1.61059e+07 muA


** Expected Voltages: 
** ibias: 1.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.83301  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.622001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 4.24801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerTransistorStack1Load2: 4.69801  V
** innerTransistorStack2Load2: 4.69801  V
** out1: 4.15001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.619001  V


.END