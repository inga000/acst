** Name: one_stage_single_output_op_amp104

.MACRO one_stage_single_output_op_amp104 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=84e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=9e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
mMainBias4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=60e-6
mTelescopicFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=428e-6
mMainBias6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=10e-6 W=10e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=84e-6
mTelescopicFirstStageLoad8 out inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=84e-6
mMainBias9 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=21e-6
mTelescopicFirstStageLoad10 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=10e-6 W=83e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=79e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=79e-6
mMainBias13 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=60e-6
mMainBias14 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=82e-6
mTelescopicFirstStageLoad15 out outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=10e-6 W=83e-6
mMainBias16 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=19e-6
mTelescopicFirstStageStageBias17 sourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=428e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp104

** Expected Performance Values: 
** Gain: 95 dB
** Power consumption: 0.547001 mW
** Area: 10965 (mu_m)^2
** Transit frequency: 3.38001 MHz
** Transit frequency with error factor: 3.37988 MHz
** Slew rate: 3.60869 V/mu_s
** Phase margin: 61.8795°
** CMRR: 147 dB
** VoutMax: 3.31001 V
** VoutMin: 0.300001 V
** VcmMax: 3.21001 V
** VcmMin: 0.610001 V


** Expected Currents: 
** NormalTransistorNmos: 8.16201e+06 muA
** NormalTransistorPmos: -3.16699e+06 muA
** NormalTransistorPmos: -1.38519e+07 muA
** NormalTransistorPmos: -3.20849e+07 muA
** NormalTransistorPmos: -3.20849e+07 muA
** DiodeTransistorNmos: 3.20841e+07 muA
** NormalTransistorNmos: 3.20841e+07 muA
** NormalTransistorNmos: 3.20841e+07 muA
** NormalTransistorPmos: -7.23299e+07 muA
** DiodeTransistorPmos: -7.23289e+07 muA
** NormalTransistorPmos: -3.20839e+07 muA
** NormalTransistorPmos: -3.20839e+07 muA
** DiodeTransistorNmos: 3.16601e+06 muA
** DiodeTransistorNmos: 1.38511e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -8.16299e+06 muA


** Expected Voltages: 
** ibias: 3.35801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.18001  V
** outVoltageBiasXXnXX0: 0.585001  V
** outVoltageBiasXXpXX2: 1.97401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.21401  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.00501  V
** sourceGCC2: 3.00501  V
** inner: 4.17701  V


.END