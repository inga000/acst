** Name: two_stage_single_output_op_amp_147_9

.MACRO two_stage_single_output_op_amp_147_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=5e-6 W=10e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mMainBias3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=7e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=541e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mMainBias6 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=19e-6
mSimpleFirstStageTransconductor7 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=25e-6
mSimpleFirstStageLoad8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=5e-6 W=8e-6
mSimpleFirstStageStageBias9 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=180e-6
mMainBias10 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=7e-6
mSecondStage1StageBias11 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=541e-6
mSimpleFirstStageLoad12 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=5e-6 W=10e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=25e-6
mSimpleFirstStageLoad14 FirstStageYinnerOutputLoad1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=225e-6
mMainBias15 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=65e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=271e-6
mSimpleFirstStageLoad17 outFirstStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=225e-6
mMainBias18 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 12.5e-12
.EOM two_stage_single_output_op_amp_147_9

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 14.9991 mW
** Area: 3997 (mu_m)^2
** Transit frequency: 8.04401 MHz
** Transit frequency with error factor: 8.03031 MHz
** Slew rate: 7.58091 V/mu_s
** Phase margin: 60.1606°
** CMRR: 88 dB
** VoutMax: 4.25 V
** VoutMin: 1.09001 V
** VcmMax: 5.23001 V
** VcmMin: 0.710001 V


** Expected Currents: 
** NormalTransistorPmos: -3.44759e+07 muA
** NormalTransistorPmos: -5.23499e+06 muA
** DiodeTransistorNmos: 7.16961e+07 muA
** DiodeTransistorNmos: 7.16951e+07 muA
** NormalTransistorNmos: 7.16941e+07 muA
** NormalTransistorNmos: 7.16951e+07 muA
** NormalTransistorPmos: -1.1931e+08 muA
** NormalTransistorPmos: -1.1931e+08 muA
** NormalTransistorNmos: 9.52311e+07 muA
** NormalTransistorNmos: 4.76161e+07 muA
** NormalTransistorNmos: 4.76161e+07 muA
** NormalTransistorNmos: 2.70157e+09 muA
** DiodeTransistorNmos: 2.70157e+09 muA
** NormalTransistorPmos: -2.70156e+09 muA
** DiodeTransistorNmos: 3.44751e+07 muA
** NormalTransistorNmos: 3.44741e+07 muA
** DiodeTransistorNmos: 5.23401e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.26401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.49401  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.747001  V
** outVoltageBiasXXnXX2: 0.563001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 2.19501  V
** innerSourceLoad1: 1.13601  V
** innerTransistorStack2Load1: 1.13701  V
** sourceTransconductance: 1.94501  V
** inner: 0.747001  V


.END