** Name: two_stage_single_output_op_amp_68_9

.MACRO two_stage_single_output_op_amp_68_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=9e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=112e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=293e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=142e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=38e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=6e-6 W=38e-6
mMainBias7 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=90e-6
mFoldedCascodeFirstStageStageBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=156e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=53e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=53e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=9e-6
mSecondStage1StageBias13 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=293e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=21e-6
mFoldedCascodeFirstStageLoad15 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=1e-6 W=38e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=44e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=44e-6
mFoldedCascodeFirstStageStageBias18 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=156e-6
mMainBias19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=90e-6
mMainBias20 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=198e-6
mMainBias21 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=599e-6
mSecondStage1Transconductor22 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=282e-6
mFoldedCascodeFirstStageLoad23 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=6e-6 W=38e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_68_9

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 4.38001 mW
** Area: 14978 (mu_m)^2
** Transit frequency: 2.93701 MHz
** Transit frequency with error factor: 2.93745 MHz
** Slew rate: 3.63319 V/mu_s
** Phase margin: 68.182°
** CMRR: 134 dB
** VoutMax: 4.25 V
** VoutMin: 1.23001 V
** VcmMax: 3.27001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.20909e+07 muA
** NormalTransistorPmos: -6.76149e+07 muA
** NormalTransistorNmos: 1.64041e+07 muA
** NormalTransistorNmos: 2.52371e+07 muA
** NormalTransistorNmos: 1.64041e+07 muA
** NormalTransistorNmos: 2.52371e+07 muA
** DiodeTransistorPmos: -1.64049e+07 muA
** NormalTransistorPmos: -1.64059e+07 muA
** NormalTransistorPmos: -1.64049e+07 muA
** DiodeTransistorPmos: -1.64059e+07 muA
** NormalTransistorPmos: -1.76639e+07 muA
** DiodeTransistorPmos: -1.76629e+07 muA
** NormalTransistorPmos: -8.83199e+06 muA
** NormalTransistorPmos: -8.83199e+06 muA
** NormalTransistorNmos: 7.15815e+08 muA
** DiodeTransistorNmos: 7.15814e+08 muA
** NormalTransistorPmos: -7.15814e+08 muA
** DiodeTransistorNmos: 2.20901e+07 muA
** NormalTransistorNmos: 2.20891e+07 muA
** DiodeTransistorNmos: 6.76141e+07 muA
** DiodeTransistorNmos: 6.76151e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.48301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.64001  V
** inputVoltageBiasXXnXX2: 1.12901  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.820001  V
** outSourceVoltageBiasXXnXX2: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.24201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.27701  V
** innerTransistorStack2Load2: 4.28001  V
** out1: 3.33401  V
** sourceGCC1: 0.531001  V
** sourceGCC2: 0.531001  V
** sourceTransconductance: 3.27501  V
** inner: 0.816001  V
** inner: 4.24001  V


.END