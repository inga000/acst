** Name: two_stage_single_output_op_amp_63_1

.MACRO two_stage_single_output_op_amp_63_1 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=5e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=86e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=4e-6 W=158e-6
m5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=8e-6
m6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m7 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=12e-6
m8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
m9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=70e-6
m10 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
m11 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=112e-6
m12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=12e-6
m13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=20e-6
m14 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=23e-6
m15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=86e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=75e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=75e-6
m18 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=8e-6 W=178e-6
m19 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=446e-6
m20 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=158e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_63_1

** Expected Performance Values: 
** Gain: 114 dB
** Power consumption: 3.61201 mW
** Area: 6448 (mu_m)^2
** Transit frequency: 3.56801 MHz
** Transit frequency with error factor: 3.56767 MHz
** Slew rate: 6.70121 V/mu_s
** Phase margin: 65.8902°
** CMRR: 135 dB
** VoutMax: 4.73001 V
** VoutMin: 0.620001 V
** VcmMax: 3.02001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.00071e+07 muA
** NormalTransistorNmos: 1.33431e+07 muA
** NormalTransistorNmos: 3.03741e+07 muA
** NormalTransistorNmos: 4.57791e+07 muA
** NormalTransistorNmos: 3.03741e+07 muA
** NormalTransistorNmos: 4.57791e+07 muA
** DiodeTransistorPmos: -3.0375e+07 muA
** DiodeTransistorPmos: -3.03759e+07 muA
** NormalTransistorPmos: -3.0375e+07 muA
** NormalTransistorPmos: -3.03759e+07 muA
** NormalTransistorPmos: -3.08129e+07 muA
** NormalTransistorPmos: -3.08139e+07 muA
** NormalTransistorPmos: -1.54059e+07 muA
** NormalTransistorPmos: -1.54059e+07 muA
** NormalTransistorNmos: 5.97517e+08 muA
** NormalTransistorPmos: -5.97516e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.00079e+07 muA
** DiodeTransistorPmos: -1.33439e+07 muA


** Expected Voltages: 
** ibias: 1.22801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 1.02301  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX2: 4.16301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.15401  V
** innerStageBias: 4.52701  V
** innerTransistorStack2Load2: 4.15301  V
** out1: 3.38201  V
** sourceGCC1: 0.522001  V
** sourceGCC2: 0.522001  V
** sourceTransconductance: 3.36601  V


.END