.suckt  symmetrical_op_amp121 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad3 out1FirstStage out1FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mSymmetricalFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad5 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mSymmetricalFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSymmetricalFirstStageTransconductor8 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1StageBias10 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
mSecondStage1StageBias11 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStage1Transconductor12 out out1FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor13 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias14 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor15 innerComplementarySecondStage inSourceTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mMainBias17 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias18 ibias ibias sourceNmos sourceNmos nmos
mMainBias19 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
.end symmetrical_op_amp121

