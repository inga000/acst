.suckt  two_stage_fully_differential_op_amp_9_3 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m5 outFeedback outFeedback sourceNmos sourceNmos nmos
m6 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m7 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m8 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m9 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m10 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m11 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m12 out1FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m13 out2FirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m14 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m15 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m16 sourceTransconductance ibias sourcePmos sourcePmos pmos
m17 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m18 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m19 out1 out1FirstStage sourceNmos sourceNmos nmos
m20 out1 inputVoltageBiasXXpXX2 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m21 SecondStage1YinnerStageBias ibias sourcePmos sourcePmos pmos
m22 out2 out2FirstStage sourceNmos sourceNmos nmos
m23 out2 inputVoltageBiasXXpXX2 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m24 SecondStage2YinnerStageBias ibias sourcePmos sourcePmos pmos
m25 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m26 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
m27 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m28 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_9_3

