** Name: two_stage_single_output_op_amp_57_1

.MACRO two_stage_single_output_op_amp_57_1 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=14e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
m3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=47e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=10e-6 W=19e-6
m5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=81e-6
m6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=22e-6
m7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=46e-6
m8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=46e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=32e-6
m10 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=22e-6
m11 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
m12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=168e-6
m13 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=15e-6
m14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=89e-6
m15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=89e-6
m16 FirstStageYsourceTransconductance outVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=10e-6 W=280e-6
m17 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=517e-6
m18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=2e-6 W=47e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_57_1

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 4.51801 mW
** Area: 5799 (mu_m)^2
** Transit frequency: 4.00901 MHz
** Transit frequency with error factor: 4.00421 MHz
** Slew rate: 4.40928 V/mu_s
** Phase margin: 69.328°
** CMRR: 102 dB
** VoutMax: 4.72001 V
** VoutMin: 0.510001 V
** VcmMax: 3.22001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.89661e+07 muA
** NormalTransistorNmos: 1.11376e+08 muA
** NormalTransistorNmos: 1.99141e+07 muA
** NormalTransistorNmos: 3.00841e+07 muA
** NormalTransistorNmos: 1.99141e+07 muA
** NormalTransistorNmos: 3.00841e+07 muA
** DiodeTransistorPmos: -1.99149e+07 muA
** NormalTransistorPmos: -1.99149e+07 muA
** NormalTransistorPmos: -2.03429e+07 muA
** NormalTransistorPmos: -2.03439e+07 muA
** NormalTransistorPmos: -1.01709e+07 muA
** NormalTransistorPmos: -1.01709e+07 muA
** NormalTransistorNmos: 7.03066e+08 muA
** NormalTransistorPmos: -7.03065e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.89669e+07 muA
** DiodeTransistorPmos: -1.11375e+08 muA


** Expected Voltages: 
** ibias: 1.12201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.917001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.16001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.45101  V
** out1: 4.21801  V
** sourceGCC1: 0.537001  V
** sourceGCC2: 0.537001  V
** sourceTransconductance: 3.24201  V


.END