** Name: two_stage_single_output_op_amp_80_7

.MACRO two_stage_single_output_op_amp_80_7 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=86e-6
mMainBias2 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=3e-6 W=96e-6
mMainBias3 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=7e-6 W=92e-6
mFoldedCascodeFirstStageStageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=12e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=4e-6 W=17e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=4e-6 W=33e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=10e-6
mFoldedCascodeFirstStageTransconductor11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=10e-6
mFoldedCascodeFirstStageStageBias12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=12e-6
mMainBias13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=92e-6
mSecondStage1StageBias14 out inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=3e-6 W=121e-6
mFoldedCascodeFirstStageLoad15 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=4e-6 W=33e-6
mFoldedCascodeFirstStageLoad16 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=40e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageLoad18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mMainBias19 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=575e-6
mMainBias20 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=446e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=10e-6 W=563e-6
mFoldedCascodeFirstStageLoad22 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=40e-6
mMainBias23 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=124e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_80_7

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 8.95201 mW
** Area: 9834 (mu_m)^2
** Transit frequency: 3.37001 MHz
** Transit frequency with error factor: 3.37006 MHz
** Slew rate: 3.58987 V/mu_s
** Phase margin: 61.3065°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.410001 V
** VcmMax: 5.17001 V
** VcmMin: 1.65001 V


** Expected Currents: 
** NormalTransistorPmos: -1.24615e+08 muA
** NormalTransistorPmos: -5.73195e+08 muA
** NormalTransistorPmos: -4.52188e+08 muA
** NormalTransistorPmos: -1.62229e+07 muA
** NormalTransistorPmos: -2.43329e+07 muA
** NormalTransistorPmos: -1.62229e+07 muA
** NormalTransistorPmos: -2.43329e+07 muA
** NormalTransistorNmos: 1.62221e+07 muA
** NormalTransistorNmos: 1.62211e+07 muA
** NormalTransistorNmos: 1.62221e+07 muA
** NormalTransistorNmos: 1.62211e+07 muA
** NormalTransistorNmos: 1.62211e+07 muA
** DiodeTransistorNmos: 1.62201e+07 muA
** NormalTransistorNmos: 8.11101e+06 muA
** NormalTransistorNmos: 8.11101e+06 muA
** NormalTransistorNmos: 5.71636e+08 muA
** NormalTransistorPmos: -5.71635e+08 muA
** DiodeTransistorNmos: 1.24616e+08 muA
** NormalTransistorNmos: 1.24615e+08 muA
** DiodeTransistorNmos: 5.73196e+08 muA
** DiodeTransistorNmos: 4.52189e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.969001  V
** inputVoltageBiasXXnXX3: 0.813001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.47601  V
** outSourceVoltageBiasXXnXX1: 0.738001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 0.411001  V
** innerTransistorStack2Load2: 0.412001  V
** out1: 0.617001  V
** sourceGCC1: 4.11201  V
** sourceGCC2: 4.11201  V
** sourceTransconductance: 1.92501  V
** inner: 0.735001  V


.END