.suckt  two_stage_single_output_op_amp_94_5 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m3 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m4 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m5 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m6 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m7 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
m8 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m9 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos
m10 sourceTransconductance ibias sourceNmos sourceNmos nmos
m11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c2 out sourceNmos 
m13 out outFirstStage sourceNmos sourceNmos nmos
m14 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m15 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m16 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
m17 ibias ibias sourceNmos sourceNmos nmos
m18 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m19 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m21 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_94_5

