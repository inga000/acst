** Name: two_stage_single_output_op_amp_45_10

.MACRO two_stage_single_output_op_amp_45_10 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=20e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=13e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=288e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=454e-6
m7 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=225e-6
m8 outVoltageBiasXXpXX1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=25e-6
m9 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=225e-6
m10 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=181e-6
m11 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=181e-6
m12 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=5e-6 W=460e-6
m13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=349e-6
m14 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=367e-6
m15 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=34e-6
m16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=288e-6
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=67e-6
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=67e-6
m19 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=507e-6
m20 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 7.40001e-12
.EOM two_stage_single_output_op_amp_45_10

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 5.04901 mW
** Area: 14954 (mu_m)^2
** Transit frequency: 3.69501 MHz
** Transit frequency with error factor: 3.69505 MHz
** Slew rate: 17.0084 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** VoutMax: 4.25 V
** VoutMin: 0.160001 V
** VcmMax: 3.47001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.63971e+07 muA
** NormalTransistorPmos: -8.72999e+07 muA
** NormalTransistorPmos: -8.44799e+06 muA
** NormalTransistorNmos: 1.28512e+08 muA
** NormalTransistorNmos: 1.92766e+08 muA
** NormalTransistorNmos: 1.28513e+08 muA
** NormalTransistorNmos: 1.92767e+08 muA
** DiodeTransistorPmos: -1.28511e+08 muA
** NormalTransistorPmos: -1.28512e+08 muA
** NormalTransistorPmos: -1.28511e+08 muA
** NormalTransistorPmos: -1.28508e+08 muA
** NormalTransistorPmos: -6.42549e+07 muA
** NormalTransistorPmos: -6.42549e+07 muA
** NormalTransistorNmos: 4.82176e+08 muA
** NormalTransistorPmos: -4.82175e+08 muA
** NormalTransistorPmos: -4.82174e+08 muA
** DiodeTransistorNmos: 8.72991e+07 muA
** DiodeTransistorNmos: 8.44701e+06 muA
** DiodeTransistorPmos: -2.63979e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.964001  V
** out: 2.5  V
** outFirstStage: 4.22501  V
** outVoltageBiasXXnXX2: 0.563001  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.56201  V
** out1: 4.27801  V
** sourceGCC1: 0.358001  V
** sourceGCC2: 0.358001  V
** sourceTransconductance: 3.79301  V
** innerTransconductance: 4.78901  V


.END