** Name: two_stage_single_output_op_amp_39_7

.MACRO two_stage_single_output_op_amp_39_7 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=11e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=62e-6
m3 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=16e-6
m4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=119e-6
m5 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=5e-6 W=119e-6
m6 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
m7 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=17e-6
m8 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=27e-6
m9 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=36e-6
m10 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=17e-6
m11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=48e-6
m12 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=171e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=358e-6
m14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=5e-6 W=119e-6
m15 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=119e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_39_7

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 4.35601 mW
** Area: 7732 (mu_m)^2
** Transit frequency: 3.71801 MHz
** Transit frequency with error factor: 3.71544 MHz
** Slew rate: 3.5037 V/mu_s
** Phase margin: 60.1606°
** CMRR: 107 dB
** negPSRR: 103 dB
** posPSRR: 98 dB
** VoutMax: 4.49001 V
** VoutMin: 0.230001 V
** VcmMax: 3.91001 V
** VcmMin: 1.34001 V


** Expected Currents: 
** NormalTransistorNmos: 2.44551e+07 muA
** NormalTransistorPmos: -2.56743e+08 muA
** DiodeTransistorPmos: -1.61909e+07 muA
** NormalTransistorPmos: -1.61919e+07 muA
** NormalTransistorPmos: -1.61909e+07 muA
** DiodeTransistorPmos: -1.61919e+07 muA
** NormalTransistorNmos: 3.23791e+07 muA
** NormalTransistorNmos: 3.23781e+07 muA
** NormalTransistorNmos: 1.61901e+07 muA
** NormalTransistorNmos: 1.61901e+07 muA
** NormalTransistorNmos: 5.47517e+08 muA
** NormalTransistorPmos: -5.47516e+08 muA
** DiodeTransistorNmos: 2.56744e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.44559e+07 muA


** Expected Voltages: 
** ibias: 0.636001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.790001  V
** out: 2.5  V
** outFirstStage: 3.92701  V
** outVoltageBiasXXpXX0: 3.85401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.26101  V
** innerStageBias: 0.231001  V
** innerTransistorStack1Load1: 4.26001  V
** out1: 3.50101  V
** sourceTransconductance: 1.94501  V


.END