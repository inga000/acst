** Name: two_stage_single_output_op_amp_65_5

.MACRO two_stage_single_output_op_amp_65_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=5e-6 W=10e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=26e-6
mMainBias3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=68e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=291e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=12e-6
mMainBias6 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=6e-6 W=88e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=16e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=78e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=78e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=105e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=16e-6
mMainBias12 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=234e-6
mMainBias13 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=63e-6
mMainBias14 outVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=42e-6
mFoldedCascodeFirstStageStageBias15 FirstStageYinnerStageBias outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=6e-6 W=111e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=74e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=74e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=206e-6
mFoldedCascodeFirstStageTransconductor19 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=61e-6
mFoldedCascodeFirstStageTransconductor20 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=61e-6
mFoldedCascodeFirstStageStageBias21 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=5e-6 W=88e-6
mMainBias22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=68e-6
mSecondStage1StageBias23 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=291e-6
mFoldedCascodeFirstStageLoad24 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=206e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.80001e-12
.EOM two_stage_single_output_op_amp_65_5

** Expected Performance Values: 
** Gain: 124 dB
** Power consumption: 2.92101 mW
** Area: 14647 (mu_m)^2
** Transit frequency: 2.80501 MHz
** Transit frequency with error factor: 2.80466 MHz
** Slew rate: 4.06834 V/mu_s
** Phase margin: 60.1606°
** CMRR: 132 dB
** VoutMax: 3 V
** VoutMin: 0.590001 V
** VcmMax: 3.14001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 8.91371e+07 muA
** NormalTransistorNmos: 2.39991e+07 muA
** NormalTransistorNmos: 1.60091e+07 muA
** NormalTransistorNmos: 1.96971e+07 muA
** NormalTransistorNmos: 2.97131e+07 muA
** NormalTransistorNmos: 1.96971e+07 muA
** NormalTransistorNmos: 2.97131e+07 muA
** NormalTransistorPmos: -1.96979e+07 muA
** NormalTransistorPmos: -1.96989e+07 muA
** NormalTransistorPmos: -1.96979e+07 muA
** NormalTransistorPmos: -1.96989e+07 muA
** NormalTransistorPmos: -2.00349e+07 muA
** NormalTransistorPmos: -2.00359e+07 muA
** NormalTransistorPmos: -1.00169e+07 muA
** NormalTransistorPmos: -1.00169e+07 muA
** NormalTransistorNmos: 3.85523e+08 muA
** NormalTransistorPmos: -3.85522e+08 muA
** DiodeTransistorPmos: -3.85523e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -8.91379e+07 muA
** NormalTransistorPmos: -8.91389e+07 muA
** DiodeTransistorPmos: -2.4e+07 muA
** DiodeTransistorPmos: -1.60099e+07 muA


** Expected Voltages: 
** ibias: 1.20201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.997001  V
** outInputVoltageBiasXXpXX1: 2.43601  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.71701  V
** outVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXpXX3: 4.18901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.50201  V
** innerTransistorStack1Load2: 4.41301  V
** innerTransistorStack2Load2: 4.41301  V
** out1: 4.04901  V
** sourceGCC1: 0.526001  V
** sourceGCC2: 0.526001  V
** sourceTransconductance: 3.29801  V
** inner: 3.71301  V


.END