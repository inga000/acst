** Name: two_stage_single_output_op_amp_50_6

.MACRO two_stage_single_output_op_amp_50_6 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYinnerLoad2 FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=267e-6
m2 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
m3 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=9e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=7e-6 W=22e-6
m5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=9e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=415e-6
m7 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=22e-6
m8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=14e-6
m9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=14e-6
m10 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=80e-6
m11 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=600e-6
m12 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
m13 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=9e-6 W=578e-6
m14 outFirstStage FirstStageYinnerLoad2 sourceNmos sourceNmos nmos4 L=4e-6 W=267e-6
m15 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=17e-6
m16 FirstStageYinnerLoad2 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=111e-6
m17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=139e-6
m18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=139e-6
m19 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=9e-6
m20 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=25e-6
m21 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=415e-6
m22 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=111e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10.5e-12
.EOM two_stage_single_output_op_amp_50_6

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 8.90301 mW
** Area: 14996 (mu_m)^2
** Transit frequency: 4.82001 MHz
** Transit frequency with error factor: 4.81757 MHz
** Slew rate: 12.139 V/mu_s
** Phase margin: 60.1606°
** CMRR: 101 dB
** VoutMax: 3 V
** VoutMin: 0.640001 V
** VcmMax: 4.66001 V
** VcmMin: 1.06001 V


** Expected Currents: 
** NormalTransistorNmos: 2.78151e+07 muA
** NormalTransistorNmos: 3.13151e+07 muA
** NormalTransistorPmos: -3.54629e+07 muA
** NormalTransistorPmos: -1.28887e+08 muA
** NormalTransistorPmos: -1.94333e+08 muA
** NormalTransistorPmos: -1.28887e+08 muA
** NormalTransistorPmos: -1.94333e+08 muA
** DiodeTransistorNmos: 1.28888e+08 muA
** NormalTransistorNmos: 1.28888e+08 muA
** NormalTransistorNmos: 1.30891e+08 muA
** NormalTransistorNmos: 6.54451e+07 muA
** NormalTransistorNmos: 6.54451e+07 muA
** NormalTransistorNmos: 1.28726e+09 muA
** NormalTransistorNmos: 1.28726e+09 muA
** NormalTransistorPmos: -1.28725e+09 muA
** DiodeTransistorPmos: -1.28725e+09 muA
** DiodeTransistorNmos: 3.54621e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.78159e+07 muA
** NormalTransistorPmos: -2.78169e+07 muA
** DiodeTransistorPmos: -3.13159e+07 muA
** DiodeTransistorPmos: -3.13169e+07 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.04901  V
** inputVoltageBiasXXpXX2: 2.37901  V
** out: 2.5  V
** outFirstStage: 0.564001  V
** outInputVoltageBiasXXpXX1: 2.43601  V
** outSourceVoltageBiasXXpXX1: 3.71801  V
** outSourceVoltageBiasXXpXX2: 3.69301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerLoad2: 0.556001  V
** sourceGCC1: 3.61501  V
** sourceGCC2: 3.61501  V
** sourceTransconductance: 1.68601  V
** innerTransconductance: 0.159001  V
** inner: 3.71701  V


.END