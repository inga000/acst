** Name: two_stage_single_output_op_amp_66_2

.MACRO two_stage_single_output_op_amp_66_2 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=9e-6 W=29e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
mMainBias3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=25e-6
mMainBias4 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=31e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=3e-6 W=311e-6
mFoldedCascodeFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=110e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=26e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC1 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=83e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC2 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=83e-6
mSecondStage1Transconductor10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=48e-6
mMainBias11 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=370e-6
mMainBias12 inputVoltageBiasXXpXX3 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=78e-6
mSecondStage1Transconductor13 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=5e-6 W=63e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=26e-6
mMainBias15 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=9e-6 W=195e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=48e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=48e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=2e-6 W=73e-6
mFoldedCascodeFirstStageTransconductor19 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=33e-6
mFoldedCascodeFirstStageTransconductor20 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=33e-6
mFoldedCascodeFirstStageStageBias21 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=110e-6
mMainBias22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=311e-6
mMainBias23 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=47e-6
mSecondStage1StageBias24 out inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=8e-6 W=151e-6
mFoldedCascodeFirstStageLoad25 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=2e-6 W=73e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.60001e-12
.EOM two_stage_single_output_op_amp_66_2

** Expected Performance Values: 
** Gain: 135 dB
** Power consumption: 2.28401 mW
** Area: 13998 (mu_m)^2
** Transit frequency: 2.56301 MHz
** Transit frequency with error factor: 2.5626 MHz
** Slew rate: 3.55725 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** VoutMax: 4.38001 V
** VoutMin: 0.530001 V
** VcmMax: 3.18001 V
** VcmMin: -0.369999 V


** Expected Currents: 
** NormalTransistorNmos: 6.62471e+07 muA
** NormalTransistorNmos: 1.26917e+08 muA
** NormalTransistorNmos: 2.64991e+07 muA
** NormalTransistorPmos: -4.08269e+07 muA
** NormalTransistorNmos: 1.64481e+07 muA
** NormalTransistorNmos: 2.81981e+07 muA
** NormalTransistorNmos: 1.64481e+07 muA
** NormalTransistorNmos: 2.81981e+07 muA
** NormalTransistorPmos: -1.64489e+07 muA
** NormalTransistorPmos: -1.64499e+07 muA
** NormalTransistorPmos: -1.64489e+07 muA
** NormalTransistorPmos: -1.64499e+07 muA
** NormalTransistorPmos: -2.34989e+07 muA
** DiodeTransistorPmos: -2.35e+07 muA
** NormalTransistorPmos: -1.17489e+07 muA
** NormalTransistorPmos: -1.17489e+07 muA
** NormalTransistorNmos: 1.2992e+08 muA
** NormalTransistorNmos: 1.29919e+08 muA
** NormalTransistorPmos: -1.29919e+08 muA
** DiodeTransistorNmos: 4.08261e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -6.62479e+07 muA
** NormalTransistorPmos: -6.62489e+07 muA
** DiodeTransistorPmos: -1.26916e+08 muA
** DiodeTransistorPmos: -2.65e+07 muA


** Expected Voltages: 
** ibias: 0.596001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.989001  V
** inputVoltageBiasXXpXX2: 3.68601  V
** inputVoltageBiasXXpXX3: 3.81501  V
** out: 2.5  V
** outFirstStage: 0.584001  V
** outInputVoltageBiasXXpXX1: 3.49201  V
** outSourceVoltageBiasXXpXX1: 4.24601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.40901  V
** innerTransistorStack2Load2: 4.40901  V
** out1: 4.04501  V
** sourceGCC1: 0.391001  V
** sourceGCC2: 0.391001  V
** sourceTransconductance: 3.37901  V
** innerTransconductance: 0.234001  V
** inner: 4.24501  V


.END