.suckt  one_stage_fully_differential_op_amp10 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
m1 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m4 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m5 outFeedback outFeedback sourceNmos sourceNmos nmos
m6 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXpXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m7 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
m8 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXpXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m9 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
m10 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m11 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m12 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m13 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m14 out1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m15 out2 outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m16 out1 outFeedback sourceNmos sourceNmos nmos
m17 out2 outFeedback sourceNmos sourceNmos nmos
m18 sourceTransconductance ibias sourcePmos sourcePmos pmos
m19 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m20 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c1 out1 sourceNmos 
c2 out2 sourceNmos 
m21 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m22 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos
m23 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m24 ibias ibias sourcePmos sourcePmos pmos
.end one_stage_fully_differential_op_amp10

