.suckt  two_stage_fully_differential_op_amp_36_4 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_3 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_4 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_5 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_Load_6 outFeedback outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_7 FeedbackStageYsourceTransconductance1 outVoltageBiasXXpXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m_FullyDifferential_FeedbackdStage_StageBias_8 FeedbackStageYinnerStageBias1 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYsourceTransconductance2 outVoltageBiasXXpXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m_FullyDifferential_FeedbackdStage_StageBias_10 FeedbackStageYinnerStageBias2 ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackStage_Transconductor_11 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m_FullyDifferential_FeedbackStage_Transconductor_13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FeedbackStage_Transconductor_14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m_FullyDifferential_FirstStage_Load_15 out1FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m_FullyDifferential_FirstStage_Load_16 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_17 out2FirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m_FullyDifferential_FirstStage_Load_18 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Load_19 out1FirstStage ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_20 out2FirstStage ibias sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_StageBias_21 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m_FullyDifferential_FirstStage_StageBias_22 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Transconductor_23 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_FullyDifferential_FirstStage_Transconductor_24 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_Transconductor_25 out1 inputVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m_FullyDifferential_SecondStage1_Transconductor_26 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_StageBias_27 out1 outVoltageBiasXXpXX2 SecondStage1YinnerStageBias SecondStage1YinnerStageBias pmos
m_FullyDifferential_SecondStage1_StageBias_28 SecondStage1YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_Transconductor_29 out2 inputVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m_FullyDifferential_SecondStage2_Transconductor_30 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_StageBias_31 out2 outVoltageBiasXXpXX2 SecondStage2YinnerStageBias SecondStage2YinnerStageBias pmos
m_FullyDifferential_SecondStage2_StageBias_32 SecondStage2YinnerStageBias ibias sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_33 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_34 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_35 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m_FullyDifferential_MainBias_36 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_37 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_38 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_36_4

