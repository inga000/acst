** Name: symmetrical_op_amp186

.MACRO symmetrical_op_amp186 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=22e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias3 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=13e-6
mSymmetricalFirstStageStageBias5 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=8e-6 W=71e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=28e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=47e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias8 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=47e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=42e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias10 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=3e-6 W=33e-6
mSecondStage1StageBias11 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=33e-6
mSymmetricalFirstStageTransconductor12 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=42e-6
mMainBias13 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=8e-6 W=112e-6
mMainBias14 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=8e-6 W=12e-6
mSymmetricalFirstStageLoad15 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=15e-6
mSymmetricalFirstStageLoad16 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=15e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=43e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=43e-6
mMainBias19 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=81e-6
mSymmetricalFirstStageLoad20 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=79e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor21 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=231e-6
mSecondStage1Transconductor22 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=231e-6
mSymmetricalFirstStageLoad23 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=79e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp186

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 1.12401 mW
** Area: 4885 (mu_m)^2
** Transit frequency: 4.85301 MHz
** Transit frequency with error factor: 4.85258 MHz
** Slew rate: 4.64389 V/mu_s
** Phase margin: 72.1927°
** CMRR: 143 dB
** negPSRR: 120 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 0.410001 V
** VcmMax: 4.81001 V
** VcmMin: 1.37001 V


** Expected Currents: 
** NormalTransistorNmos: 5.38701e+06 muA
** NormalTransistorNmos: 5.07661e+07 muA
** NormalTransistorPmos: -3.35379e+07 muA
** NormalTransistorPmos: -1.6e+07 muA
** NormalTransistorPmos: -1.60009e+07 muA
** NormalTransistorPmos: -1.6e+07 muA
** NormalTransistorPmos: -1.60009e+07 muA
** NormalTransistorNmos: 3.19971e+07 muA
** NormalTransistorNmos: 3.19961e+07 muA
** NormalTransistorNmos: 1.59991e+07 muA
** NormalTransistorNmos: 1.59991e+07 muA
** NormalTransistorNmos: 4.65701e+07 muA
** NormalTransistorNmos: 4.65691e+07 muA
** NormalTransistorPmos: -4.65709e+07 muA
** NormalTransistorPmos: -4.65699e+07 muA
** NormalTransistorNmos: 4.65701e+07 muA
** NormalTransistorNmos: 4.65691e+07 muA
** NormalTransistorPmos: -4.65709e+07 muA
** NormalTransistorPmos: -4.65699e+07 muA
** DiodeTransistorNmos: 3.35371e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.38799e+06 muA
** DiodeTransistorPmos: -5.07669e+07 muA


** Expected Voltages: 
** ibias: 0.612001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.815001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.592001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 4.22001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.208001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.187001  V
** innerTransconductance: 4.40001  V
** inner: 0.187001  V
** inner: 4.40001  V


.END