.suckt  symmetrical_op_amp114 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos
mMainBias2 out2FirstStage ibias sourceNmos sourceNmos nmos
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad4 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
mSymmetricalFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageLoad6 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
mSymmetricalFirstStageLoad7 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mSymmetricalFirstStageStageBias8 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
mSymmetricalFirstStageTransconductor9 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
mSymmetricalFirstStageTransconductor10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
cLoadCapacitor1 out sourceNmos 
mSecondStage1StageBias11 out outVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos
mSecondStage1StageBias12 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStage1Transconductor13 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
mSecondStage1Transconductor14 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
mSecondStageWithVoltageBiasAsStageBiasStageBias15 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos
mSecondStageWithVoltageBiasAsStageBiasTransconductor17 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos
mMainBias18 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
mMainBias19 ibias ibias sourceNmos sourceNmos nmos
mMainBias20 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
mMainBias21 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos
.end symmetrical_op_amp114

