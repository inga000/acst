** Name: two_stage_single_output_op_amp_45_1

.MACRO two_stage_single_output_op_amp_45_1 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=7e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
m3 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
m4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=7e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=194e-6
m6 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=65e-6
m7 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=10e-6
m8 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
m9 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=31e-6
m10 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=10e-6
m11 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
m12 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
m13 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=313e-6
m14 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=4e-6 W=32e-6
m15 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=194e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=150e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=9e-6 W=150e-6
m18 FirstStageYsourceTransconductance outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_45_1

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 5.01301 mW
** Area: 6086 (mu_m)^2
** Transit frequency: 3.62201 MHz
** Transit frequency with error factor: 3.62185 MHz
** Slew rate: 3.84143 V/mu_s
** Phase margin: 73.9116°
** CMRR: 142 dB
** VoutMax: 4.43001 V
** VoutMin: 0.580001 V
** VcmMax: 3.69001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.26761e+07 muA
** NormalTransistorNmos: 2.06691e+07 muA
** NormalTransistorNmos: 1.73221e+07 muA
** NormalTransistorNmos: 2.61601e+07 muA
** NormalTransistorNmos: 1.73221e+07 muA
** NormalTransistorNmos: 2.61601e+07 muA
** DiodeTransistorPmos: -1.73229e+07 muA
** NormalTransistorPmos: -1.73229e+07 muA
** NormalTransistorPmos: -1.73229e+07 muA
** NormalTransistorPmos: -1.76789e+07 muA
** NormalTransistorPmos: -8.83899e+06 muA
** NormalTransistorPmos: -8.83899e+06 muA
** NormalTransistorNmos: 9.06862e+08 muA
** NormalTransistorPmos: -9.06861e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.26769e+07 muA
** DiodeTransistorPmos: -2.06699e+07 muA


** Expected Voltages: 
** ibias: 1.18701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.982001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 3.86401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.59701  V
** out1: 4.27801  V
** sourceGCC1: 0.533001  V
** sourceGCC2: 0.533001  V
** sourceTransconductance: 3.23601  V


.END