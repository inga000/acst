** Name: two_stage_single_output_op_amp_167_3

.MACRO two_stage_single_output_op_amp_167_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=239e-6
mSimpleFirstStageLoad2 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=154e-6
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=4e-6 W=478e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=24e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mSimpleFirstStageLoad6 FirstStageYout1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=324e-6
mSecondStage1Transconductor7 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=496e-6
mSimpleFirstStageLoad8 outFirstStage outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=324e-6
mSimpleFirstStageStageBias9 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
mSimpleFirstStageLoad10 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=154e-6
mSimpleFirstStageTransconductor11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=77e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=45e-6
mSecondStage1StageBias13 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=311e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=598e-6
mSimpleFirstStageLoad15 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=478e-6
mSimpleFirstStageTransconductor16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=77e-6
mMainBias17 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=291e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 6.5e-12
.EOM two_stage_single_output_op_amp_167_3

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 7.16001 mW
** Area: 12757 (mu_m)^2
** Transit frequency: 4.39401 MHz
** Transit frequency with error factor: 4.35206 MHz
** Slew rate: 5.58358 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.03001 V
** VoutMin: 0.150001 V
** VcmMax: 3.22001 V
** VcmMin: -0.289999 V


** Expected Currents: 
** NormalTransistorPmos: -2.92053e+08 muA
** DiodeTransistorPmos: -3.8357e+08 muA
** DiodeTransistorPmos: -3.83571e+08 muA
** NormalTransistorPmos: -3.8357e+08 muA
** NormalTransistorPmos: -3.83571e+08 muA
** NormalTransistorNmos: 4.02328e+08 muA
** NormalTransistorNmos: 4.02328e+08 muA
** NormalTransistorPmos: -3.75139e+07 muA
** NormalTransistorPmos: -3.75129e+07 muA
** NormalTransistorPmos: -1.87569e+07 muA
** NormalTransistorPmos: -1.87569e+07 muA
** NormalTransistorNmos: 3.15317e+08 muA
** NormalTransistorPmos: -3.15316e+08 muA
** NormalTransistorPmos: -3.15315e+08 muA
** DiodeTransistorNmos: 2.92054e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.48201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.675001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.68601  V
** innerStageBias: 4.26101  V
** innerTransistorStack2Load1: 3.68301  V
** out1: 2.69701  V
** sourceTransconductance: 3.26601  V
** innerStageBias: 4.21701  V


.END