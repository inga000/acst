** Name: symmetrical_op_amp55

.MACRO symmetrical_op_amp55 ibias in1 in2 out sourceNmos sourcePmos
m1 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=21e-6
m2 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=10e-6 W=11e-6
m3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=21e-6
m4 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=61e-6
m5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=41e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=131e-6
m7 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=10e-6 W=12e-6
m8 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=10e-6 W=12e-6
m9 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=46e-6
m10 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=46e-6
m11 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=37e-6
m12 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=215e-6
m13 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=61e-6
m14 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=2e-6 W=8e-6
m15 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=37e-6
m16 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=131e-6
m17 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=41e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp55

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 0.876001 mW
** Area: 3566 (mu_m)^2
** Transit frequency: 3.60601 MHz
** Transit frequency with error factor: 3.60563 MHz
** Slew rate: 3.50002 V/mu_s
** Phase margin: 78.4953°
** CMRR: 141 dB
** negPSRR: 44 dB
** posPSRR: 45 dB
** VoutMax: 3.37001 V
** VoutMin: 0.75 V
** VcmMax: 3.25 V
** VcmMin: 0.0100001 V


** Expected Currents: 
** NormalTransistorPmos: -5.29069e+07 muA
** DiodeTransistorNmos: 1.61841e+07 muA
** DiodeTransistorNmos: 1.61841e+07 muA
** NormalTransistorPmos: -3.23699e+07 muA
** DiodeTransistorPmos: -3.23689e+07 muA
** NormalTransistorPmos: -1.61849e+07 muA
** NormalTransistorPmos: -1.61849e+07 muA
** NormalTransistorNmos: 3.50071e+07 muA
** NormalTransistorNmos: 3.50061e+07 muA
** NormalTransistorPmos: -3.50079e+07 muA
** DiodeTransistorPmos: -3.50089e+07 muA
** NormalTransistorPmos: -3.49899e+07 muA
** NormalTransistorNmos: 3.49891e+07 muA
** NormalTransistorNmos: 3.49881e+07 muA
** DiodeTransistorNmos: 5.29061e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40201  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 1.15501  V
** inSourceTransconductanceComplementarySecondStage: 0.570001  V
** inStageBiasComplementarySecondStage: 4.07601  V
** innerComplementarySecondStage: 2.80901  V
** out: 2.5  V
** outFirstStage: 0.570001  V
** outSourceVoltageBiasXXpXX1: 4.20201  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.22001  V
** innerTransconductance: 0.165001  V
** inner: 0.165001  V
** inner: 4.19901  V


.END