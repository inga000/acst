** Name: one_stage_single_output_op_amp81

.MACRO one_stage_single_output_op_amp81 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=7e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=85e-6
m4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=9e-6 W=85e-6
m5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=19e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=16e-6
m7 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=41e-6
m8 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=9e-6 W=85e-6
m9 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=116e-6
m10 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=85e-6
m11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=40e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=40e-6
m13 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=115e-6
m14 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=362e-6
m15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=362e-6
m16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=65e-6
m17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=65e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp81

** Expected Performance Values: 
** Gain: 87 dB
** Power consumption: 1.30201 mW
** Area: 4860 (mu_m)^2
** Transit frequency: 4.02001 MHz
** Transit frequency with error factor: 4.02008 MHz
** Slew rate: 3.65578 V/mu_s
** Phase margin: 84.7978°
** CMRR: 142 dB
** VoutMax: 3.85001 V
** VoutMin: 0.880001 V
** VcmMax: 4.97001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 2.71621e+07 muA
** NormalTransistorPmos: -7.35099e+07 muA
** NormalTransistorPmos: -1.11603e+08 muA
** NormalTransistorPmos: -7.35099e+07 muA
** NormalTransistorPmos: -1.11603e+08 muA
** DiodeTransistorNmos: 7.35091e+07 muA
** NormalTransistorNmos: 7.35081e+07 muA
** NormalTransistorNmos: 7.35091e+07 muA
** DiodeTransistorNmos: 7.35081e+07 muA
** NormalTransistorNmos: 7.61851e+07 muA
** NormalTransistorNmos: 7.61841e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.71629e+07 muA
** DiodeTransistorPmos: -2.71639e+07 muA


** Expected Voltages: 
** ibias: 1.18701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 3.99801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.580001  V
** innerStageBias: 0.629001  V
** innerTransistorStack1Load2: 0.578001  V
** out1: 1.28701  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.94501  V


.END