** Name: two_stage_single_output_op_amp_68_3

.MACRO two_stage_single_output_op_amp_68_3 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=9e-6 W=33e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=47e-6
m3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=16e-6
m4 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=3e-6 W=4e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=127e-6
m6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=4e-6
m7 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=62e-6
m8 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=10e-6 W=62e-6
m9 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=9e-6 W=42e-6
m10 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=177e-6
m11 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=10e-6
m12 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=41e-6
m13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=9e-6 W=42e-6
m14 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=119e-6
m15 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=119e-6
m16 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=10e-6 W=62e-6
m17 out outInputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=3e-6 W=167e-6
m18 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=62e-6
m19 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=88e-6
m20 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=88e-6
m21 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=127e-6
m22 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=243e-6
m23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=16e-6
Capacitor1 outFirstStage out 4.5e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_68_3

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 2.95101 mW
** Area: 11359 (mu_m)^2
** Transit frequency: 2.86101 MHz
** Transit frequency with error factor: 2.86113 MHz
** Slew rate: 3.70188 V/mu_s
** Phase margin: 61.3065°
** CMRR: 133 dB
** VoutMax: 3.12001 V
** VoutMin: 0.530001 V
** VcmMax: 3.24001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 2.11901e+06 muA
** NormalTransistorNmos: 8.69101e+06 muA
** NormalTransistorNmos: 1.67601e+07 muA
** NormalTransistorNmos: 2.51841e+07 muA
** NormalTransistorNmos: 1.67601e+07 muA
** NormalTransistorNmos: 2.51841e+07 muA
** DiodeTransistorPmos: -1.67609e+07 muA
** NormalTransistorPmos: -1.67619e+07 muA
** NormalTransistorPmos: -1.67609e+07 muA
** DiodeTransistorPmos: -1.67619e+07 muA
** NormalTransistorPmos: -1.68509e+07 muA
** DiodeTransistorPmos: -1.68519e+07 muA
** NormalTransistorPmos: -8.42499e+06 muA
** NormalTransistorPmos: -8.42499e+06 muA
** NormalTransistorNmos: 5.18921e+08 muA
** NormalTransistorPmos: -5.1892e+08 muA
** NormalTransistorPmos: -5.18921e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.11999e+06 muA
** NormalTransistorPmos: -2.12099e+06 muA
** DiodeTransistorPmos: -8.69199e+06 muA
** DiodeTransistorPmos: -8.69299e+06 muA


** Expected Voltages: 
** ibias: 1.13901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.934001  V
** outInputVoltageBiasXXpXX1: 3.44801  V
** outInputVoltageBiasXXpXX2: 2.66401  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.22401  V
** outSourceVoltageBiasXXpXX2: 3.83501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.26201  V
** innerTransistorStack1Load2: 4.25901  V
** out1: 3.30801  V
** sourceGCC1: 0.527001  V
** sourceGCC2: 0.527001  V
** sourceTransconductance: 3.27001  V
** innerStageBias: 3.94701  V
** inner: 4.22201  V


.END