.suckt  symmetrical_op_amp13 ibias in1 in2 out sourceNmos sourcePmos
m1 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos
m2 outFirstStage outFirstStage sourceNmos sourceNmos nmos
m3 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m4 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m5 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m6 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c1 out sourceNmos 
m7 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m9 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos
m10 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m11 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos
m12 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m13 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m14 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m15 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp13

