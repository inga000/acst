** Name: two_stage_single_output_op_amp_47_10

.MACRO two_stage_single_output_op_amp_47_10 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=62e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=34e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=33e-6
m4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=48e-6
m5 out inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=552e-6
m6 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=158e-6
m7 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=255e-6
m8 FirstStageYinnerSourceLoad2 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=158e-6
m9 FirstStageYsourceGCC1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=107e-6
m10 FirstStageYsourceGCC2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=1e-6 W=107e-6
m11 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
m12 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=391e-6
m13 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=93e-6
m14 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=479e-6
m15 FirstStageYinnerSourceLoad2 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=93e-6
m16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=384e-6
m17 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=384e-6
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=41e-6
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=41e-6
m20 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=556e-6
m21 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=344e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 19.2001e-12
.EOM two_stage_single_output_op_amp_47_10

** Expected Performance Values: 
** Gain: 126 dB
** Power consumption: 11.1651 mW
** Area: 12165 (mu_m)^2
** Transit frequency: 4.13601 MHz
** Transit frequency with error factor: 4.1361 MHz
** Slew rate: 6.21294 V/mu_s
** Phase margin: 60.1606°
** CMRR: 134 dB
** VoutMax: 4.27001 V
** VoutMin: 0.150001 V
** VcmMax: 3.84001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 4.87363e+08 muA
** NormalTransistorPmos: -1.46063e+08 muA
** NormalTransistorPmos: -1.18087e+08 muA
** NormalTransistorNmos: 1.19642e+08 muA
** NormalTransistorNmos: 2.05101e+08 muA
** NormalTransistorNmos: 1.19638e+08 muA
** NormalTransistorNmos: 2.05095e+08 muA
** NormalTransistorPmos: -1.19639e+08 muA
** NormalTransistorPmos: -1.19638e+08 muA
** NormalTransistorPmos: -1.19637e+08 muA
** NormalTransistorPmos: -1.19638e+08 muA
** NormalTransistorPmos: -1.70915e+08 muA
** NormalTransistorPmos: -8.54579e+07 muA
** NormalTransistorPmos: -8.54579e+07 muA
** NormalTransistorNmos: 1.05136e+09 muA
** NormalTransistorPmos: -1.05135e+09 muA
** NormalTransistorPmos: -1.05135e+09 muA
** DiodeTransistorNmos: 1.46064e+08 muA
** DiodeTransistorNmos: 1.18088e+08 muA
** DiodeTransistorPmos: -4.87362e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.17501  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.555001  V
** out: 2.5  V
** outFirstStage: 4.02101  V
** outVoltageBiasXXnXX1: 1.00401  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.24901  V
** innerTransistorStack1Load2: 4.51701  V
** innerTransistorStack2Load2: 4.51701  V
** sourceGCC1: 0.350001  V
** sourceGCC2: 0.350001  V
** sourceTransconductance: 3.40401  V
** innerTransconductance: 4.56201  V


.END