.suckt  two_stage_fully_differential_op_amp_24_2 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXpXX1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m2 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 inputVoltageBiasXXnXX3 ibias sourcePmos sourcePmos pmos
m5 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m6 outFeedback outFeedback sourcePmos sourcePmos pmos
m7 FeedbackStageYsourceTransconductance1 inputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m8 FeedbackStageYinnerStageBias1 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m9 FeedbackStageYsourceTransconductance2 inputVoltageBiasXXnXX2 FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m10 FeedbackStageYinnerStageBias2 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m11 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m12 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m13 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m14 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m15 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m16 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m17 out1FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos
m18 FirstStageYinnerTransistorStack1Load2 outFeedback sourcePmos sourcePmos pmos
m19 out2FirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos
m20 FirstStageYinnerTransistorStack2Load2 outFeedback sourcePmos sourcePmos pmos
m21 sourceTransconductance inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m22 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m23 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m24 out1 inputVoltageBiasXXnXX2 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m25 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m26 out1 ibias sourcePmos sourcePmos pmos
m27 out2 inputVoltageBiasXXnXX2 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m28 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m29 out2 ibias sourcePmos sourcePmos pmos
m30 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
m31 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m32 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m33 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m34 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_24_2

