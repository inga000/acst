.suckt  two_stage_fully_differential_op_amp_17_1 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m4 outFeedback outFeedback sourcePmos sourcePmos pmos
m5 FeedbackStageYsourceTransconductance1 ibias sourceNmos sourceNmos nmos
m6 FeedbackStageYsourceTransconductance2 ibias sourceNmos sourceNmos nmos
m7 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m8 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m9 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m10 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m11 out1FirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m12 FirstStageYsourceGCC1 outFeedback sourcePmos sourcePmos pmos
m13 out2FirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m14 FirstStageYsourceGCC2 outFeedback sourcePmos sourcePmos pmos
m15 out1FirstStage ibias sourceNmos sourceNmos nmos
m16 out2FirstStage ibias sourceNmos sourceNmos nmos
m17 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m20 out1 out1FirstStage sourceNmos sourceNmos nmos
m21 out1 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m22 out2 out2FirstStage sourceNmos sourceNmos nmos
m23 out2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m24 ibias ibias sourceNmos sourceNmos nmos
m25 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m26 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_17_1

