** Name: symmetrical_op_amp97

.MACRO symmetrical_op_amp97 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=22e-6
mMainBias2 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=37e-6
mSecondStage1StageBias3 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=160e-6
mSymmetricalFirstStageLoad4 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=41e-6
mSymmetricalFirstStageLoad5 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=41e-6
mSecondStage1Transconductor6 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=52e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor7 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=52e-6
mSymmetricalFirstStageLoad8 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=30e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=2e-6 W=38e-6
mSecondStage1Transconductor10 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=38e-6
mSymmetricalFirstStageLoad11 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=30e-6
mSymmetricalFirstStageStageBias12 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=571e-6
mSymmetricalFirstStageTransconductor13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=105e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias14 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=160e-6
mSecondStage1StageBias15 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=2e-6 W=130e-6
mSymmetricalFirstStageTransconductor16 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=105e-6
mMainBias17 out2FirstStage ibias sourcePmos sourcePmos pmos4 L=4e-6 W=537e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp97

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 2.60901 mW
** Area: 5872 (mu_m)^2
** Transit frequency: 7.73801 MHz
** Transit frequency with error factor: 7.73769 MHz
** Slew rate: 9.9379 V/mu_s
** Phase margin: 86.5167°
** CMRR: 147 dB
** negPSRR: 48 dB
** posPSRR: 159 dB
** VoutMax: 3.96001 V
** VoutMin: 0.400001 V
** VcmMax: 3.99001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.46038e+08 muA
** NormalTransistorNmos: 7.86001e+07 muA
** NormalTransistorNmos: 7.85991e+07 muA
** NormalTransistorNmos: 7.86001e+07 muA
** NormalTransistorNmos: 7.85991e+07 muA
** NormalTransistorPmos: -1.57201e+08 muA
** NormalTransistorPmos: -7.86009e+07 muA
** NormalTransistorPmos: -7.86009e+07 muA
** NormalTransistorNmos: 9.95611e+07 muA
** NormalTransistorNmos: 9.95601e+07 muA
** NormalTransistorPmos: -9.95619e+07 muA
** DiodeTransistorPmos: -9.95629e+07 muA
** NormalTransistorPmos: -9.90409e+07 muA
** NormalTransistorNmos: 9.90401e+07 muA
** NormalTransistorNmos: 9.90411e+07 muA
** DiodeTransistorNmos: 1.46039e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18901  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** inStageBiasComplementarySecondStage: 4.24901  V
** innerComplementarySecondStage: 3.39101  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.803001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.26801  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END