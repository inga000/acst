.suckt  symmetrical_op_amp89 ibias in1 in2 out sourceNmos sourcePmos
m_Symmetrical_FirstStage_Load_1 out2FirstStage out2FirstStage out1FirstStage out1FirstStage nmos
m_Symmetrical_FirstStage_Load_2 out1FirstStage out1FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_Load_3 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage nmos
m_Symmetrical_FirstStage_Load_4 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_FirstStage_StageBias_5 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m_Symmetrical_FirstStage_Transconductor_6 out2FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_Symmetrical_FirstStage_Transconductor_7 inOutputTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_Symmetrical_Load_Capacitor_1 out sourceNmos 
m_Symmetrical_SecondStage1_Transconductor_8 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m_Symmetrical_SecondStage1_Transconductor_9 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m_Symmetrical_SecondStage1_StageBias_10 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m_Symmetrical_SecondStage1_StageBias_11 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_12 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_StageBias_13 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_14 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m_Symmetrical_SecondStageWithVoltageBiasAsStageBias_Transconductor_15 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m_Symmetrical_MainBias_16 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp89

