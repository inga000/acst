** Name: two_stage_single_output_op_amp_81_7

.MACRO two_stage_single_output_op_amp_81_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=48e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=48e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=49e-6
mMainBias5 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=10e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=17e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=48e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=14e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=14e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=10e-6
mSecondStage1StageBias12 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=6e-6 W=384e-6
mFoldedCascodeFirstStageLoad13 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=48e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=46e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=28e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=10e-6 W=429e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=46e-6
mMainBias19 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=434e-6
mMainBias20 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=55e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_81_7

** Expected Performance Values: 
** Gain: 117 dB
** Power consumption: 5.03801 mW
** Area: 9074 (mu_m)^2
** Transit frequency: 2.51601 MHz
** Transit frequency with error factor: 2.51549 MHz
** Slew rate: 4.12999 V/mu_s
** Phase margin: 61.8795°
** CMRR: 144 dB
** VoutMax: 4.25 V
** VoutMin: 0.280001 V
** VcmMax: 5.17001 V
** VcmMin: 1.52001 V


** Expected Currents: 
** NormalTransistorPmos: -4.40022e+08 muA
** NormalTransistorPmos: -5.52079e+07 muA
** NormalTransistorPmos: -1.86819e+07 muA
** NormalTransistorPmos: -2.83879e+07 muA
** NormalTransistorPmos: -1.86819e+07 muA
** NormalTransistorPmos: -2.83879e+07 muA
** DiodeTransistorNmos: 1.86811e+07 muA
** NormalTransistorNmos: 1.86801e+07 muA
** NormalTransistorNmos: 1.86811e+07 muA
** DiodeTransistorNmos: 1.86801e+07 muA
** NormalTransistorNmos: 1.94091e+07 muA
** NormalTransistorNmos: 1.94081e+07 muA
** NormalTransistorNmos: 9.70501e+06 muA
** NormalTransistorNmos: 9.70501e+06 muA
** NormalTransistorNmos: 4.35581e+08 muA
** NormalTransistorPmos: -4.3558e+08 muA
** DiodeTransistorNmos: 4.40023e+08 muA
** DiodeTransistorNmos: 5.52071e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.39801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 1.04001  V
** outVoltageBiasXXnXX2: 0.689001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.484001  V
** innerTransistorStack1Load2: 0.583001  V
** innerTransistorStack2Load2: 0.584001  V
** out1: 1.14001  V
** sourceGCC1: 4.11201  V
** sourceGCC2: 4.11201  V
** sourceTransconductance: 1.82301  V


.END