** Name: two_stage_single_output_op_amp_68_3

.MACRO two_stage_single_output_op_amp_68_3 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=7e-6 W=17e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mFoldedCascodeFirstStageLoad3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=102e-6
mFoldedCascodeFirstStageLoad4 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=10e-6 W=102e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=7e-6 W=66e-6
mMainBias6 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=205e-6
mMainBias8 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=24e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=100e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=100e-6
mSecondStage1Transconductor12 out outFirstStage sourceNmos sourceNmos nmos4 L=6e-6 W=201e-6
mFoldedCascodeFirstStageLoad13 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=24e-6
mMainBias14 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=22e-6
mMainBias15 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=88e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=3e-6 W=102e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=146e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=146e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=205e-6
mSecondStage1StageBias20 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=372e-6
mMainBias21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=66e-6
mSecondStage1StageBias22 out outInputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=188e-6
mFoldedCascodeFirstStageLoad23 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=10e-6 W=102e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_68_3

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 5.05301 mW
** Area: 13445 (mu_m)^2
** Transit frequency: 3.85101 MHz
** Transit frequency with error factor: 3.85074 MHz
** Slew rate: 3.99904 V/mu_s
** Phase margin: 67.6091°
** CMRR: 137 dB
** VoutMax: 3.54001 V
** VoutMin: 0.570001 V
** VcmMax: 3.33001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 6.00601e+06 muA
** NormalTransistorNmos: 2.45091e+07 muA
** NormalTransistorNmos: 1.81041e+07 muA
** NormalTransistorNmos: 2.73001e+07 muA
** NormalTransistorNmos: 1.81041e+07 muA
** NormalTransistorNmos: 2.73001e+07 muA
** DiodeTransistorPmos: -1.81049e+07 muA
** NormalTransistorPmos: -1.81059e+07 muA
** NormalTransistorPmos: -1.81049e+07 muA
** DiodeTransistorPmos: -1.81059e+07 muA
** NormalTransistorPmos: -1.83949e+07 muA
** DiodeTransistorPmos: -1.83959e+07 muA
** NormalTransistorPmos: -9.19699e+06 muA
** NormalTransistorPmos: -9.19699e+06 muA
** NormalTransistorNmos: 9.15426e+08 muA
** NormalTransistorPmos: -9.15425e+08 muA
** NormalTransistorPmos: -9.15426e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -6.00699e+06 muA
** NormalTransistorPmos: -6.00799e+06 muA
** DiodeTransistorPmos: -2.45099e+07 muA
** DiodeTransistorPmos: -2.45109e+07 muA


** Expected Voltages: 
** ibias: 1.18101  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.976001  V
** outInputVoltageBiasXXpXX1: 3.49601  V
** outInputVoltageBiasXXpXX2: 3.12801  V
** outSourceVoltageBiasXXnXX1: 0.556001  V
** outSourceVoltageBiasXXpXX1: 4.24801  V
** outSourceVoltageBiasXXpXX2: 4.06401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.26101  V
** innerTransistorStack2Load2: 4.26301  V
** out1: 3.38301  V
** sourceGCC1: 0.525001  V
** sourceGCC2: 0.525001  V
** sourceTransconductance: 3.23201  V
** innerStageBias: 4.21201  V
** inner: 4.24801  V


.END