** Name: two_stage_single_output_op_amp_43_9

.MACRO two_stage_single_output_op_amp_43_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=62e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=6e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=294e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=56e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=82e-6
m6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=11e-6
m7 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=294e-6
m8 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=36e-6
m9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=36e-6
m10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=48e-6
m11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=48e-6
m12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
m13 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=263e-6
m14 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=485e-6
m15 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=11e-6
m16 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=107e-6
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=141e-6
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=141e-6
m19 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=281e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 6.80001e-12
.EOM two_stage_single_output_op_amp_43_9

** Expected Performance Values: 
** Gain: 83 dB
** Power consumption: 4.26201 mW
** Area: 13276 (mu_m)^2
** Transit frequency: 3.43501 MHz
** Transit frequency with error factor: 3.42691 MHz
** Slew rate: 5.03454 V/mu_s
** Phase margin: 60.1606°
** CMRR: 89 dB
** VoutMax: 4.25 V
** VoutMin: 1.20001 V
** VcmMax: 4 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorPmos: -1.31459e+07 muA
** NormalTransistorPmos: -5.93279e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 5.14251e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 5.14251e+07 muA
** DiodeTransistorPmos: -3.42849e+07 muA
** NormalTransistorPmos: -3.42849e+07 muA
** NormalTransistorPmos: -3.42849e+07 muA
** NormalTransistorPmos: -1.71419e+07 muA
** NormalTransistorPmos: -1.71419e+07 muA
** NormalTransistorNmos: 6.5702e+08 muA
** DiodeTransistorNmos: 6.57019e+08 muA
** NormalTransistorPmos: -6.57019e+08 muA
** DiodeTransistorNmos: 1.31451e+07 muA
** NormalTransistorNmos: 1.31441e+07 muA
** DiodeTransistorNmos: 5.93271e+07 muA
** DiodeTransistorNmos: 5.93281e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.23301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.11901  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.60201  V
** outSourceVoltageBiasXXnXX1: 0.801001  V
** outSourceVoltageBiasXXnXX2: 0.564001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.71001  V
** sourceGCC1: 0.564001  V
** sourceGCC2: 0.564001  V
** sourceTransconductance: 3.29701  V
** inner: 0.801001  V


.END