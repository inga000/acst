** Name: two_stage_single_output_op_amp_189_9

.MACRO two_stage_single_output_op_amp_189_9 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=32e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=6e-6 W=6e-6
mMainBias3 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=8e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=83e-6
mMainBias5 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=5e-6 W=63e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=10e-6
mSimpleFirstStageStageBias8 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=13e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=28e-6
mSimpleFirstStageLoad10 FirstStageYout1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=9e-6 W=32e-6
mSimpleFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=21e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSecondStage1StageBias13 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=6e-6 W=83e-6
mSimpleFirstStageLoad14 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=6e-6 W=42e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=28e-6
mSimpleFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=174e-6
mSimpleFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=174e-6
mSimpleFirstStageLoad18 FirstStageYout1 ibias FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=5e-6 W=600e-6
mMainBias19 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=42e-6
mMainBias20 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=10e-6
mSecondStage1Transconductor21 out outFirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=233e-6
mSimpleFirstStageLoad22 outFirstStage ibias FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=600e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_189_9

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 5.09201 mW
** Area: 12096 (mu_m)^2
** Transit frequency: 3.15601 MHz
** Transit frequency with error factor: 3.15357 MHz
** Slew rate: 3.90533 V/mu_s
** Phase margin: 61.8795°
** CMRR: 120 dB
** VoutMax: 4.25 V
** VoutMin: 1.82001 V
** VcmMax: 4.59001 V
** VcmMin: 1.62001 V


** Expected Currents: 
** NormalTransistorPmos: -4.27519e+07 muA
** NormalTransistorPmos: -9.97799e+06 muA
** NormalTransistorNmos: 1.67924e+08 muA
** NormalTransistorNmos: 1.67925e+08 muA
** DiodeTransistorNmos: 1.67924e+08 muA
** NormalTransistorPmos: -1.77115e+08 muA
** NormalTransistorPmos: -1.77114e+08 muA
** NormalTransistorPmos: -1.77115e+08 muA
** NormalTransistorPmos: -1.77114e+08 muA
** NormalTransistorNmos: 1.83831e+07 muA
** NormalTransistorNmos: 1.83821e+07 muA
** NormalTransistorNmos: 9.19201e+06 muA
** NormalTransistorNmos: 9.19201e+06 muA
** NormalTransistorNmos: 5.91436e+08 muA
** DiodeTransistorNmos: 5.91435e+08 muA
** NormalTransistorPmos: -5.91435e+08 muA
** DiodeTransistorNmos: 4.27511e+07 muA
** NormalTransistorNmos: 4.27501e+07 muA
** DiodeTransistorNmos: 9.97701e+06 muA
** DiodeTransistorNmos: 9.97601e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 2.22601  V
** inputVoltageBiasXXnXX2: 1.47201  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 1.11301  V
** outSourceVoltageBiasXXnXX2: 0.747001  V
** outSourceVoltageBiasXXpXX1: 3.90501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15501  V
** innerStageBias: 0.797001  V
** innerTransistorStack1Load2: 3.98001  V
** innerTransistorStack2Load2: 3.98001  V
** out1: 2.09501  V
** sourceTransconductance: 1.89801  V
** inner: 1.10701  V


.END