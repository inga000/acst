** Name: two_stage_single_output_op_amp_61_1

.MACRO two_stage_single_output_op_amp_61_1 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=7e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=88e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=5e-6 W=17e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=15e-6
mFoldedCascodeFirstStageLoad7 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=64e-6
mFoldedCascodeFirstStageLoad8 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=64e-6
mMainBias9 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=52e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=105e-6
mFoldedCascodeFirstStageLoad11 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=15e-6
mMainBias12 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mFoldedCascodeFirstStageStageBias13 FirstStageYinnerStageBias outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=20e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=88e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=16e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=16e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=5e-6 W=347e-6
mSecondStage1StageBias18 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=2e-6 W=525e-6
mFoldedCascodeFirstStageLoad19 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=5e-6 W=325e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_61_1

** Expected Performance Values: 
** Gain: 116 dB
** Power consumption: 4.34601 mW
** Area: 7174 (mu_m)^2
** Transit frequency: 3.11701 MHz
** Transit frequency with error factor: 3.1174 MHz
** Slew rate: 6.11517 V/mu_s
** Phase margin: 73.3387°
** CMRR: 131 dB
** VoutMax: 4.60001 V
** VoutMin: 0.580001 V
** VcmMax: 3.01001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 3.45201e+07 muA
** NormalTransistorNmos: 8.53301e+06 muA
** NormalTransistorNmos: 2.78951e+07 muA
** NormalTransistorNmos: 4.18551e+07 muA
** NormalTransistorNmos: 2.78951e+07 muA
** NormalTransistorNmos: 4.18551e+07 muA
** DiodeTransistorPmos: -2.78959e+07 muA
** NormalTransistorPmos: -2.78959e+07 muA
** NormalTransistorPmos: -2.78959e+07 muA
** NormalTransistorPmos: -2.79229e+07 muA
** NormalTransistorPmos: -2.79239e+07 muA
** NormalTransistorPmos: -1.39609e+07 muA
** NormalTransistorPmos: -1.39609e+07 muA
** NormalTransistorNmos: 7.32466e+08 muA
** NormalTransistorPmos: -7.32465e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -3.45209e+07 muA
** DiodeTransistorPmos: -8.53399e+06 muA


** Expected Voltages: 
** ibias: 1.18701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 0.982001  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXpXX2: 4.03901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.40001  V
** innerTransistorStack2Load2: 4.40501  V
** out1: 4.05801  V
** sourceGCC1: 0.524001  V
** sourceGCC2: 0.524001  V
** sourceTransconductance: 3.375  V


.END