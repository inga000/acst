** Name: two_stage_single_output_op_amp_53_1

.MACRO two_stage_single_output_op_amp_53_1 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=35e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=6e-6 W=50e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=26e-6
mMainBias5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=31e-6
mFoldedCascodeFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=35e-6
mFoldedCascodeFirstStageTransconductor7 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=30e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=30e-6
mFoldedCascodeFirstStageStageBias9 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=10e-6 W=135e-6
mSecondStage1Transconductor10 out outFirstStage sourceNmos sourceNmos nmos4 L=10e-6 W=299e-6
mFoldedCascodeFirstStageLoad11 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=6e-6 W=50e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=459e-6
mMainBias13 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=209e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=38e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
mSecondStage1StageBias17 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=596e-6
mFoldedCascodeFirstStageLoad18 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=38e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_53_1

** Expected Performance Values: 
** Gain: 118 dB
** Power consumption: 4.77401 mW
** Area: 14081 (mu_m)^2
** Transit frequency: 4.23501 MHz
** Transit frequency with error factor: 4.23508 MHz
** Slew rate: 3.97589 V/mu_s
** Phase margin: 64.1713°
** CMRR: 139 dB
** VoutMax: 4.73001 V
** VoutMin: 0.550001 V
** VcmMax: 5.14001 V
** VcmMin: 0.770001 V


** Expected Currents: 
** NormalTransistorNmos: 8.79951e+07 muA
** NormalTransistorNmos: 3.98891e+07 muA
** NormalTransistorPmos: -1.79979e+07 muA
** NormalTransistorPmos: -3.08549e+07 muA
** NormalTransistorPmos: -1.79959e+07 muA
** NormalTransistorPmos: -3.08529e+07 muA
** DiodeTransistorNmos: 1.79971e+07 muA
** DiodeTransistorNmos: 1.79961e+07 muA
** NormalTransistorNmos: 1.79951e+07 muA
** NormalTransistorNmos: 1.79961e+07 muA
** NormalTransistorNmos: 2.57131e+07 muA
** NormalTransistorNmos: 1.28561e+07 muA
** NormalTransistorNmos: 1.28561e+07 muA
** NormalTransistorNmos: 7.55305e+08 muA
** NormalTransistorPmos: -7.55304e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -8.79959e+07 muA
** DiodeTransistorPmos: -3.98899e+07 muA


** Expected Voltages: 
** ibias: 0.555001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.954001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.16901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.595001  V
** innerTransistorStack2Load2: 0.594001  V
** out1: 1.15901  V
** sourceGCC1: 4.53101  V
** sourceGCC2: 4.53101  V
** sourceTransconductance: 1.88101  V


.END