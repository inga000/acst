.suckt  complementary_op_amp5 ibias in1 in2 out sourceNmos sourcePmos
m_Complementary_MainBias_1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_Complementary_MainBias_2 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_3 FirstStageYinnerOutputLoadPmos outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1LoadNmos FirstStageYinnerTransistorStack1LoadNmos nmos
m_Complementary_FirstStage_Load_4 FirstStageYinnerTransistorStack1LoadNmos outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_5 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m_Complementary_FirstStage_Load_6 FirstStageYinnerTransistorStack2LoadNmos outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_7 FirstStageYinnerOutputLoadPmos FirstStageYinnerOutputLoadPmos FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos pmos
m_Complementary_FirstStage_Load_8 FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_9 out FirstStageYinnerOutputLoadPmos FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m_Complementary_FirstStage_Load_10 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_StageBias_11 FirstStageYsourceTransconductanceNmos outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_12 FirstStageYsourceTransconductancePmos ibias sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Transconductor_13 FirstStageYinnerSourceLoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_14 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_15 FirstStageYinnerTransistorStack1LoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m_Complementary_FirstStage_Transconductor_16 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c_Complementary_Load_Capacitor_1 out sourceNmos 
m_Complementary_MainBias_17 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_MainBias_18 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_Complementary_MainBias_19 ibias ibias sourcePmos sourcePmos pmos
.end complementary_op_amp5

