** Name: one_stage_single_output_op_amp115

.MACRO one_stage_single_output_op_amp115 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=15e-6
mMainBias2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos4 L=6e-6 W=8e-6
mTelescopicFirstStageLoad4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=15e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=7e-6
mTelescopicFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=135e-6
mTelescopicFirstStageLoad7 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=6e-6 W=123e-6
mTelescopicFirstStageTransconductor8 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=62e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=62e-6
mTelescopicFirstStageLoad10 out outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=6e-6 W=123e-6
mMainBias11 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=11e-6
mTelescopicFirstStageStageBias12 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=140e-6
mTelescopicFirstStageLoad13 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=15e-6
mTelescopicFirstStageLoad14 out FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=96e-6
mMainBias15 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=10e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp115

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 0.531001 mW
** Area: 3162 (mu_m)^2
** Transit frequency: 4.16101 MHz
** Transit frequency with error factor: 4.16144 MHz
** Slew rate: 4.42812 V/mu_s
** Phase margin: 80.7871°
** CMRR: 156 dB
** VoutMax: 3.51001 V
** VoutMin: 0.600001 V
** VcmMax: 3.77001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 7.23001e+06 muA
** NormalTransistorPmos: -1.01569e+07 muA
** NormalTransistorNmos: 3.93631e+07 muA
** NormalTransistorNmos: 3.93621e+07 muA
** NormalTransistorPmos: -3.93639e+07 muA
** NormalTransistorPmos: -3.93629e+07 muA
** DiodeTransistorPmos: -3.93639e+07 muA
** NormalTransistorNmos: 8.88831e+07 muA
** NormalTransistorNmos: 8.88821e+07 muA
** NormalTransistorNmos: 3.93631e+07 muA
** NormalTransistorNmos: 3.93631e+07 muA
** DiodeTransistorNmos: 1.01561e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -7.23099e+06 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX2: 0.558001  V
** outVoltageBiasXXnXX1: 2.65001  V
** outVoltageBiasXXpXX0: 3.85001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerSourceLoad2: 3.66601  V
** innerStageBias: 0.561001  V
** out1: 2.95001  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V


.END