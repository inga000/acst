** Name: symmetrical_op_amp154

.MACRO symmetrical_op_amp154 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=4e-6 W=24e-6
m2 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=1e-6 W=110e-6
m3 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=38e-6
m4 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=110e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=599e-6
m6 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=4e-6 W=54e-6
m7 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=4e-6 W=59e-6
m8 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=59e-6
m9 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=4e-6 W=54e-6
m10 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=83e-6
m11 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=83e-6
m12 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=91e-6
m13 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=2e-6 W=91e-6
m14 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=155e-6
m15 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=110e-6
m16 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=155e-6
m17 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=335e-6
m18 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=599e-6
m19 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=110e-6
m20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=38e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp154

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 2.20501 mW
** Area: 8882 (mu_m)^2
** Transit frequency: 8.18901 MHz
** Transit frequency with error factor: 8.18885 MHz
** Slew rate: 8.70347 V/mu_s
** Phase margin: 77.9223°
** CMRR: 150 dB
** negPSRR: 49 dB
** posPSRR: 161 dB
** VoutMax: 4.01001 V
** VoutMin: 0.410001 V
** VcmMax: 3.22001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -8.75079e+07 muA
** NormalTransistorNmos: 7.98061e+07 muA
** NormalTransistorNmos: 7.98051e+07 muA
** NormalTransistorNmos: 7.98061e+07 muA
** NormalTransistorNmos: 7.98051e+07 muA
** NormalTransistorPmos: -1.59613e+08 muA
** DiodeTransistorPmos: -1.59612e+08 muA
** NormalTransistorPmos: -7.98069e+07 muA
** NormalTransistorPmos: -7.98069e+07 muA
** NormalTransistorNmos: 8.71961e+07 muA
** NormalTransistorNmos: 8.71951e+07 muA
** NormalTransistorPmos: -8.71969e+07 muA
** DiodeTransistorPmos: -8.71979e+07 muA
** DiodeTransistorPmos: -8.66609e+07 muA
** NormalTransistorPmos: -8.66619e+07 muA
** NormalTransistorNmos: 8.66601e+07 muA
** NormalTransistorNmos: 8.66611e+07 muA
** DiodeTransistorNmos: 8.75071e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.38401  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 4.22501  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** innerComplementarySecondStage: 3.45001  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.818001  V
** outSourceVoltageBiasXXpXX1: 4.19301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.150001  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.23301  V
** innerTransconductance: 0.150001  V
** inner: 4.22301  V
** inner: 0.150001  V
** inner: 4.19001  V


.END