.suckt  two_stage_single_output_op_amp_199_1 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_2 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_3 FirstStageYinnerSourceLoad1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m_SingleOutput_FirstStage_Load_4 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_5 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m_SingleOutput_FirstStage_Load_6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_7 FirstStageYinnerSourceLoad1 ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_8 outFirstStage ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_StageBias_9 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos
m_SingleOutput_FirstStage_StageBias_10 FirstStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Transconductor_11 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m_SingleOutput_FirstStage_Transconductor_12 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_Transconductor_13 out outFirstStage sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_14 out ibias sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_15 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_16 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_17 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_199_1

