** Name: two_stage_single_output_op_amp_58_9

.MACRO two_stage_single_output_op_amp_58_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=8e-6 W=135e-6
m2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=21e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=148e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=109e-6
m5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=10e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=26e-6
m7 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=15e-6
m8 out inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=148e-6
m9 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=8e-6 W=41e-6
m10 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=8e-6 W=41e-6
m11 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=66e-6
m12 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=66e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=21e-6
m14 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=51e-6
m15 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=274e-6
m16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=193e-6
m17 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=15e-6
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=131e-6
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=131e-6
m20 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=26e-6
m21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 5.10001e-12
.EOM two_stage_single_output_op_amp_58_9

** Expected Performance Values: 
** Gain: 90 dB
** Power consumption: 11.6781 mW
** Area: 6277 (mu_m)^2
** Transit frequency: 5.48301 MHz
** Transit frequency with error factor: 5.47983 MHz
** Slew rate: 3.62772 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** VoutMax: 4.25 V
** VoutMin: 1.19001 V
** VcmMax: 3.05001 V
** VcmMin: -0.349999 V


** Expected Currents: 
** NormalTransistorPmos: -2.74515e+08 muA
** NormalTransistorPmos: -5.18089e+07 muA
** NormalTransistorNmos: 1.85441e+07 muA
** NormalTransistorNmos: 3.17911e+07 muA
** NormalTransistorNmos: 1.85421e+07 muA
** NormalTransistorNmos: 3.17871e+07 muA
** DiodeTransistorPmos: -1.85429e+07 muA
** NormalTransistorPmos: -1.85429e+07 muA
** NormalTransistorPmos: -2.64919e+07 muA
** DiodeTransistorPmos: -2.64909e+07 muA
** NormalTransistorPmos: -1.32459e+07 muA
** NormalTransistorPmos: -1.32459e+07 muA
** NormalTransistorNmos: 1.92566e+09 muA
** DiodeTransistorNmos: 1.92566e+09 muA
** NormalTransistorPmos: -1.92565e+09 muA
** DiodeTransistorNmos: 2.74516e+08 muA
** NormalTransistorNmos: 2.74515e+08 muA
** DiodeTransistorNmos: 5.18081e+07 muA
** DiodeTransistorNmos: 5.18091e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.19701  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.59201  V
** inputVoltageBiasXXnXX2: 1.21301  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.796001  V
** outSourceVoltageBiasXXnXX2: 0.618001  V
** outSourceVoltageBiasXXpXX1: 4.10001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 3.68901  V
** sourceGCC1: 0.601001  V
** sourceGCC2: 0.601001  V
** sourceTransconductance: 3.21401  V
** inner: 0.793001  V
** inner: 4.09401  V


.END