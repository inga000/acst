** Name: two_stage_single_output_op_amp_33_10

.MACRO two_stage_single_output_op_amp_33_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=9e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
m3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
m4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=52e-6
m5 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=305e-6
m6 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
m7 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=183e-6
m8 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=42e-6
m9 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=50e-6
m10 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=42e-6
m11 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=368e-6
m12 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=1e-6 W=211e-6
m13 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
m14 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=499e-6
m15 outVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=8e-6 W=160e-6
m16 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=2e-6 W=305e-6
m17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=333e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 19.5e-12
.EOM two_stage_single_output_op_amp_33_10

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 7.51101 mW
** Area: 11481 (mu_m)^2
** Transit frequency: 4.32901 MHz
** Transit frequency with error factor: 4.31819 MHz
** Slew rate: 16.7822 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** negPSRR: 99 dB
** posPSRR: 90 dB
** VoutMax: 4.42001 V
** VoutMin: 0.25 V
** VcmMax: 4.42001 V
** VcmMin: 1.96001 V


** Expected Currents: 
** NormalTransistorNmos: 5.45711e+07 muA
** NormalTransistorNmos: 2.03068e+08 muA
** NormalTransistorPmos: -1.64967e+08 muA
** DiodeTransistorPmos: -2.01211e+08 muA
** NormalTransistorPmos: -2.01211e+08 muA
** NormalTransistorPmos: -2.01211e+08 muA
** NormalTransistorNmos: 4.02422e+08 muA
** NormalTransistorNmos: 4.02421e+08 muA
** NormalTransistorNmos: 2.01212e+08 muA
** NormalTransistorNmos: 2.01212e+08 muA
** NormalTransistorNmos: 6.67195e+08 muA
** NormalTransistorPmos: -6.67194e+08 muA
** NormalTransistorPmos: -6.67195e+08 muA
** DiodeTransistorNmos: 1.64968e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -5.45719e+07 muA
** DiodeTransistorPmos: -2.03067e+08 muA


** Expected Voltages: 
** ibias: 0.660001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.10201  V
** outVoltageBiasXXnXX1: 0.810001  V
** outVoltageBiasXXpXX0: 3.75401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.16301  V
** innerStageBias: 0.255001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.34501  V
** innerTransconductance: 4.49901  V


.END