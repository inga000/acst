** Name: two_stage_single_output_op_amp_62_9

.MACRO two_stage_single_output_op_amp_62_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=5e-6 W=7e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=25e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=480e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=18e-6
mFoldedCascodeFirstStageLoad5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=162e-6
mMainBias6 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=6e-6 W=78e-6
mFoldedCascodeFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=274e-6
mMainBias8 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=39e-6
mFoldedCascodeFirstStageLoad9 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=25e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=117e-6
mFoldedCascodeFirstStageLoad11 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=117e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=25e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=480e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=25e-6
mMainBias15 outVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=597e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=162e-6
mFoldedCascodeFirstStageTransconductor17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=28e-6
mFoldedCascodeFirstStageTransconductor18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=28e-6
mFoldedCascodeFirstStageStageBias19 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=6e-6 W=274e-6
mMainBias20 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=78e-6
mMainBias21 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=63e-6
mSecondStage1Transconductor22 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=182e-6
mFoldedCascodeFirstStageLoad23 outFirstStage outVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=87e-6
mMainBias24 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=6e-6 W=370e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 7.10001e-12
.EOM two_stage_single_output_op_amp_62_9

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 6.89901 mW
** Area: 14204 (mu_m)^2
** Transit frequency: 4.21801 MHz
** Transit frequency with error factor: 4.21801 MHz
** Slew rate: 5.00311 V/mu_s
** Phase margin: 60.1606°
** CMRR: 139 dB
** VoutMax: 4.25 V
** VoutMin: 0.700001 V
** VcmMax: 3.27001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorNmos: 2.73462e+08 muA
** NormalTransistorPmos: -4.77369e+07 muA
** NormalTransistorPmos: -8.11799e+06 muA
** NormalTransistorNmos: 3.56651e+07 muA
** NormalTransistorNmos: 5.34961e+07 muA
** NormalTransistorNmos: 3.56661e+07 muA
** NormalTransistorNmos: 5.34971e+07 muA
** DiodeTransistorPmos: -3.56659e+07 muA
** NormalTransistorPmos: -3.56669e+07 muA
** NormalTransistorPmos: -3.56659e+07 muA
** NormalTransistorPmos: -3.56629e+07 muA
** DiodeTransistorPmos: -3.56619e+07 muA
** NormalTransistorPmos: -1.78319e+07 muA
** NormalTransistorPmos: -1.78319e+07 muA
** NormalTransistorNmos: 9.23455e+08 muA
** DiodeTransistorNmos: 9.23454e+08 muA
** NormalTransistorPmos: -9.23454e+08 muA
** DiodeTransistorNmos: 4.77361e+07 muA
** NormalTransistorNmos: 4.77351e+07 muA
** DiodeTransistorNmos: 8.11701e+06 muA
** DiodeTransistorNmos: 8.11601e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -2.73461e+08 muA


** Expected Voltages: 
** ibias: 3.45401  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.23501  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.569001  V
** outSourceVoltageBiasXXpXX1: 4.22801  V
** outVoltageBiasXXpXX2: 3.80701  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 4.52201  V
** out1: 4.21301  V
** sourceGCC1: 0.539001  V
** sourceGCC2: 0.539001  V
** sourceTransconductance: 3.25201  V
** inner: 0.555001  V
** inner: 4.22501  V


.END