** Name: two_stage_single_output_op_amp_114_8

.MACRO two_stage_single_output_op_amp_114_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=7e-6 W=12e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=10e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=17e-6
mMainBias4 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
mMainBias5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=4e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=151e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=7e-6
mTelescopicFirstStageLoad8 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=3e-6 W=24e-6
mTelescopicFirstStageTransconductor9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=40e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=40e-6
mSecondStage1StageBias11 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=7e-6 W=600e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=10e-6
mMainBias13 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=7e-6 W=15e-6
mSecondStage1StageBias14 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=7e-6 W=153e-6
mTelescopicFirstStageLoad15 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=3e-6 W=24e-6
mTelescopicFirstStageStageBias16 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=17e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=391e-6
mTelescopicFirstStageLoad18 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=4e-6 W=151e-6
mMainBias19 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=40e-6
mMainBias20 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=17e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 9.5e-12
.EOM two_stage_single_output_op_amp_114_8

** Expected Performance Values: 
** Gain: 106 dB
** Power consumption: 1.22801 mW
** Area: 8369 (mu_m)^2
** Transit frequency: 3.38701 MHz
** Transit frequency with error factor: 3.38471 MHz
** Slew rate: 4.24554 V/mu_s
** Phase margin: 60.1606°
** CMRR: 106 dB
** VoutMax: 4.85001 V
** VoutMin: 0.860001 V
** VcmMax: 4.54001 V
** VcmMin: 1.29001 V


** Expected Currents: 
** NormalTransistorNmos: 4.09501e+06 muA
** NormalTransistorPmos: -2.38479e+07 muA
** NormalTransistorPmos: -1.00589e+07 muA
** NormalTransistorNmos: 1.52381e+07 muA
** NormalTransistorNmos: 1.52381e+07 muA
** DiodeTransistorPmos: -1.52389e+07 muA
** NormalTransistorPmos: -1.52389e+07 muA
** NormalTransistorNmos: 4.05331e+07 muA
** DiodeTransistorNmos: 4.05321e+07 muA
** NormalTransistorNmos: 1.52381e+07 muA
** NormalTransistorNmos: 1.52381e+07 muA
** NormalTransistorNmos: 1.6711e+08 muA
** NormalTransistorNmos: 1.67109e+08 muA
** NormalTransistorPmos: -1.67109e+08 muA
** DiodeTransistorNmos: 2.38471e+07 muA
** NormalTransistorNmos: 2.38461e+07 muA
** DiodeTransistorNmos: 1.00581e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -4.09599e+06 muA


** Expected Voltages: 
** ibias: 1.22301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.95501  V
** out: 2.5  V
** outFirstStage: 4.28101  V
** outInputVoltageBiasXXnXX1: 1.14401  V
** outSourceVoltageBiasXXnXX1: 0.572001  V
** outSourceVoltageBiasXXnXX3: 0.556001  V
** outVoltageBiasXXnXX2: 2.65001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.28501  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerStageBias: 0.518001  V
** inner: 0.571001  V


.END