** Name: two_stage_single_output_op_amp_53_10

.MACRO two_stage_single_output_op_amp_53_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=5e-6
m2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=20e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=8e-6 W=13e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=100e-6
m5 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=132e-6
m6 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=406e-6
m7 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=172e-6
m8 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=8e-6 W=13e-6
m9 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=25e-6
m10 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=8e-6 W=20e-6
m11 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=85e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=85e-6
m13 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=36e-6
m14 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=3e-6 W=590e-6
m15 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=411e-6
m16 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=411e-6
m17 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=289e-6
m18 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=7e-6 W=289e-6
m19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=600e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 12.6001e-12
.EOM two_stage_single_output_op_amp_53_10

** Expected Performance Values: 
** Gain: 130 dB
** Power consumption: 7.08301 mW
** Area: 14266 (mu_m)^2
** Transit frequency: 3.98401 MHz
** Transit frequency with error factor: 3.98411 MHz
** Slew rate: 5.54591 V/mu_s
** Phase margin: 60.1606°
** CMRR: 128 dB
** VoutMax: 4.25 V
** VoutMin: 0.260001 V
** VcmMax: 5.03001 V
** VcmMin: 0.890001 V


** Expected Currents: 
** NormalTransistorNmos: 3.38446e+08 muA
** NormalTransistorNmos: 4.90481e+07 muA
** NormalTransistorPmos: -7.06289e+07 muA
** NormalTransistorPmos: -1.05941e+08 muA
** NormalTransistorPmos: -7.06329e+07 muA
** NormalTransistorPmos: -1.05947e+08 muA
** DiodeTransistorNmos: 7.06301e+07 muA
** DiodeTransistorNmos: 7.06311e+07 muA
** NormalTransistorNmos: 7.06321e+07 muA
** NormalTransistorNmos: 7.06311e+07 muA
** NormalTransistorNmos: 7.06291e+07 muA
** NormalTransistorNmos: 3.53141e+07 muA
** NormalTransistorNmos: 3.53141e+07 muA
** NormalTransistorNmos: 8.07172e+08 muA
** NormalTransistorPmos: -8.07171e+08 muA
** NormalTransistorPmos: -8.0717e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.38445e+08 muA
** DiodeTransistorPmos: -4.90489e+07 muA


** Expected Voltages: 
** ibias: 0.670001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.16301  V
** outVoltageBiasXXpXX2: 4.05601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.980001  V
** innerTransistorStack2Load2: 0.973001  V
** out1: 2.09801  V
** sourceGCC1: 4.41901  V
** sourceGCC2: 4.42001  V
** sourceTransconductance: 1.87301  V
** innerTransconductance: 4.72701  V


.END