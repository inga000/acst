.suckt  two_stage_single_output_op_amp_127_10 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_2 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_3 FirstStageYinnerLoad1 FirstStageYinnerLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_4 outFirstStage FirstStageYinnerLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYinnerLoad1 ibias sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_6 outFirstStage ibias sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_StageBias_7 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Transconductor_8 FirstStageYinnerLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_SingleOutput_FirstStage_Transconductor_9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_StageBias_10 out ibias sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_Transconductor_11 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos
m_SingleOutput_SecondStage1_Transconductor_12 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_13 ibias ibias sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_14 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_15 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_127_10

