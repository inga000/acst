.suckt  two_stage_fully_differential_op_amp_5_2 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m2 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m3 outFeedback outFeedback sourceNmos sourceNmos nmos
m4 FeedbackStageYsourceTransconductance1 ibias sourcePmos sourcePmos pmos
m5 FeedbackStageYsourceTransconductance2 ibias sourcePmos sourcePmos pmos
m6 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m7 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m8 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m9 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m10 out1FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m11 FirstStageYsourceGCC1 outFeedback sourceNmos sourceNmos nmos
m12 out2FirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m13 FirstStageYsourceGCC2 outFeedback sourceNmos sourceNmos nmos
m14 out1FirstStage ibias sourcePmos sourcePmos pmos
m15 out2FirstStage ibias sourcePmos sourcePmos pmos
m16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m17 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m18 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m19 out1 outVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m20 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m21 out1 ibias sourcePmos sourcePmos pmos
m22 out2 outVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m23 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m24 out2 ibias sourcePmos sourcePmos pmos
m25 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m26 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_5_2

