** Name: two_stage_single_output_op_amp_74_3

.MACRO two_stage_single_output_op_amp_74_3 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=6e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=135e-6
m3 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=403e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=52e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=268e-6
m6 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=1e-6 W=35e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=358e-6
m8 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=319e-6
m9 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=5e-6 W=403e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
m11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=8e-6
m12 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=135e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
m14 outFirstStage outInputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=265e-6
m15 out outInputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=342e-6
m16 FirstStageYout1 outInputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=265e-6
m17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=135e-6
m18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=135e-6
m19 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=562e-6
Capacitor1 outFirstStage out 10.6001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_74_3

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 10.9091 mW
** Area: 11146 (mu_m)^2
** Transit frequency: 5.77201 MHz
** Transit frequency with error factor: 5.77163 MHz
** Slew rate: 14.4979 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** VoutMax: 3.68001 V
** VoutMin: 0.580001 V
** VcmMax: 5.07001 V
** VcmMin: 1.86001 V


** Expected Currents: 
** NormalTransistorNmos: 5.27977e+08 muA
** NormalTransistorPmos: -1.54612e+08 muA
** NormalTransistorPmos: -2.65051e+08 muA
** NormalTransistorPmos: -1.54611e+08 muA
** NormalTransistorPmos: -2.6505e+08 muA
** NormalTransistorNmos: 1.54613e+08 muA
** NormalTransistorNmos: 1.54612e+08 muA
** DiodeTransistorNmos: 1.54613e+08 muA
** NormalTransistorNmos: 2.20877e+08 muA
** DiodeTransistorNmos: 2.20878e+08 muA
** NormalTransistorNmos: 1.10439e+08 muA
** NormalTransistorNmos: 1.10439e+08 muA
** NormalTransistorNmos: 1.11379e+09 muA
** NormalTransistorPmos: -1.11378e+09 muA
** NormalTransistorPmos: -1.11378e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -5.27976e+08 muA
** DiodeTransistorPmos: -5.27977e+08 muA


** Expected Voltages: 
** ibias: 1.29201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.983001  V
** outInputVoltageBiasXXpXX1: 2.78901  V
** outSourceVoltageBiasXXnXX1: 0.647001  V
** outSourceVoltageBiasXXpXX1: 4.10301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** out1: 1.18801  V
** sourceGCC1: 3.53301  V
** sourceGCC2: 3.53301  V
** sourceTransconductance: 1.52201  V
** innerStageBias: 3.77801  V
** inner: 0.643001  V


.END