** Name: two_stage_single_output_op_amp_55_3

.MACRO two_stage_single_output_op_amp_55_3 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
m2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=20e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=20e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=65e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=125e-6
m6 out outFirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=139e-6
m7 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=336e-6
m8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=20e-6
m9 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=2e-6 W=20e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=10e-6
m11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=10e-6
m12 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=7e-6 W=91e-6
m13 out inputVoltageBiasXXpXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=7e-6 W=567e-6
m14 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=27e-6
m15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=27e-6
m16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=43e-6
m17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=43e-6
m18 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=567e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_55_3

** Expected Performance Values: 
** Gain: 117 dB
** Power consumption: 2.91201 mW
** Area: 14762 (mu_m)^2
** Transit frequency: 2.51101 MHz
** Transit frequency with error factor: 2.51081 MHz
** Slew rate: 3.87689 V/mu_s
** Phase margin: 60.1606°
** CMRR: 131 dB
** VoutMax: 3.36001 V
** VoutMin: 0.5 V
** VcmMax: 4.87001 V
** VcmMin: 0.880001 V


** Expected Currents: 
** NormalTransistorNmos: 9.32961e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -3.14699e+07 muA
** NormalTransistorPmos: -1.90479e+07 muA
** NormalTransistorPmos: -3.14699e+07 muA
** DiodeTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 1.90471e+07 muA
** DiodeTransistorNmos: 1.90471e+07 muA
** NormalTransistorNmos: 2.48431e+07 muA
** NormalTransistorNmos: 1.24211e+07 muA
** NormalTransistorNmos: 1.24211e+07 muA
** NormalTransistorNmos: 4.16068e+08 muA
** NormalTransistorPmos: -4.16067e+08 muA
** NormalTransistorPmos: -4.16068e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -9.32969e+07 muA
** DiodeTransistorPmos: -9.32959e+07 muA


** Expected Voltages: 
** ibias: 0.556001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 2.58401  V
** out: 2.5  V
** outFirstStage: 0.905001  V
** outSourceVoltageBiasXXpXX1: 3.89801  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.555001  V
** innerTransistorStack1Load2: 0.555001  V
** out1: 1.11001  V
** sourceGCC1: 3.67201  V
** sourceGCC2: 3.67201  V
** sourceTransconductance: 1.77301  V
** innerStageBias: 3.68201  V


.END