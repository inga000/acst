** Name: symmetrical_op_amp185

.MACRO symmetrical_op_amp185 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=10e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=116e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=3e-6 W=27e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias5 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=14e-6
mSymmetricalFirstStageStageBias6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=83e-6
mSymmetricalFirstStageStageBias7 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=82e-6
mSecondStage1StageBias8 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=116e-6
mSymmetricalFirstStageTransconductor9 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=86e-6
mSecondStage1StageBias10 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=3e-6 W=15e-6
mSymmetricalFirstStageTransconductor11 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=86e-6
mMainBias12 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=143e-6
mSymmetricalFirstStageLoad13 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
mSymmetricalFirstStageLoad14 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
mSecondStage1Transconductor15 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=54e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor16 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=3e-6 W=54e-6
mSymmetricalFirstStageLoad17 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=101e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=289e-6
mSecondStage1Transconductor19 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=289e-6
mSymmetricalFirstStageLoad20 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=101e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp185

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 2.34001 mW
** Area: 3398 (mu_m)^2
** Transit frequency: 12.3091 MHz
** Transit frequency with error factor: 12.3088 MHz
** Slew rate: 11.6589 V/mu_s
** Phase margin: 77.9223°
** CMRR: 139 dB
** negPSRR: 128 dB
** posPSRR: 65 dB
** VoutMax: 4.25 V
** VoutMin: 1.12001 V
** VcmMax: 4.81001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorNmos: 1.42147e+08 muA
** NormalTransistorPmos: -4.09509e+07 muA
** NormalTransistorPmos: -4.09519e+07 muA
** NormalTransistorPmos: -4.09509e+07 muA
** NormalTransistorPmos: -4.09519e+07 muA
** NormalTransistorNmos: 8.18991e+07 muA
** NormalTransistorNmos: 8.18981e+07 muA
** NormalTransistorNmos: 4.09501e+07 muA
** NormalTransistorNmos: 4.09501e+07 muA
** NormalTransistorNmos: 1.16968e+08 muA
** NormalTransistorNmos: 1.16967e+08 muA
** NormalTransistorPmos: -1.16967e+08 muA
** NormalTransistorPmos: -1.16966e+08 muA
** DiodeTransistorNmos: 1.16966e+08 muA
** DiodeTransistorNmos: 1.16965e+08 muA
** NormalTransistorPmos: -1.16965e+08 muA
** NormalTransistorPmos: -1.16966e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.42146e+08 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 0.594001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 1.38901  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.557001  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.456001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V


.END