** Name: two_stage_single_output_op_amp_57_7

.MACRO two_stage_single_output_op_amp_57_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=47e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=434e-6
m3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m5 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
m7 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=89e-6
m8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=89e-6
m9 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=53e-6
m10 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=53e-6
m11 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=314e-6
m12 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
m13 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=270e-6
m14 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=541e-6
m15 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=49e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=206e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=206e-6
m18 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=27e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.80001e-12
.EOM two_stage_single_output_op_amp_57_7

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 8.70101 mW
** Area: 8440 (mu_m)^2
** Transit frequency: 3.46501 MHz
** Transit frequency with error factor: 3.45956 MHz
** Slew rate: 4.31477 V/mu_s
** Phase margin: 60.1606°
** CMRR: 90 dB
** VoutMax: 4.36001 V
** VoutMin: 0.170001 V
** VcmMax: 3.08001 V
** VcmMin: -0.389999 V


** Expected Currents: 
** NormalTransistorPmos: -2.73746e+08 muA
** NormalTransistorPmos: -5.44325e+08 muA
** NormalTransistorNmos: 4.23781e+07 muA
** NormalTransistorNmos: 6.72181e+07 muA
** NormalTransistorNmos: 4.23781e+07 muA
** NormalTransistorNmos: 6.72181e+07 muA
** DiodeTransistorPmos: -4.23789e+07 muA
** NormalTransistorPmos: -4.23789e+07 muA
** NormalTransistorPmos: -4.96809e+07 muA
** NormalTransistorPmos: -4.96799e+07 muA
** NormalTransistorPmos: -2.48409e+07 muA
** NormalTransistorPmos: -2.48409e+07 muA
** NormalTransistorNmos: 7.67725e+08 muA
** NormalTransistorPmos: -7.67724e+08 muA
** DiodeTransistorNmos: 2.73747e+08 muA
** DiodeTransistorNmos: 5.44326e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.79301  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.928001  V
** outVoltageBiasXXnXX2: 0.578001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.29301  V
** out1: 3.82201  V
** sourceGCC1: 0.373001  V
** sourceGCC2: 0.373001  V
** sourceTransconductance: 3.29601  V


.END