** Name: symmetrical_op_amp192

.MACRO symmetrical_op_amp192 ibias in1 in2 out sourceNmos sourcePmos
m1 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=9e-6 W=108e-6
m2 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=10e-6
m3 innerComplementarySecondStage innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage nmos4 L=9e-6 W=21e-6
m4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=78e-6
m5 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
m6 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=17e-6
m7 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=9e-6 W=103e-6
m8 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=17e-6
m9 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=25e-6
m10 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=78e-6
m11 SecondStageYinnerStageBias inSourceStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=9e-6 W=108e-6
m12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
m13 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=190e-6
m14 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=215e-6
m15 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=215e-6
m16 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=190e-6
m17 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=36e-6
m18 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=36e-6
m19 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=6e-6 W=40e-6
m20 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=6e-6 W=40e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp192

** Expected Performance Values: 
** Gain: 97 dB
** Power consumption: 0.994001 mW
** Area: 6474 (mu_m)^2
** Transit frequency: 2.93201 MHz
** Transit frequency with error factor: 2.93188 MHz
** Slew rate: 4.31651 V/mu_s
** Phase margin: 82.506°
** CMRR: 140 dB
** negPSRR: 115 dB
** posPSRR: 62 dB
** VoutMax: 4.25 V
** VoutMin: 0.820001 V
** VcmMax: 4.81001 V
** VcmMin: 1.47001 V


** Expected Currents: 
** NormalTransistorNmos: 2.51641e+07 muA
** NormalTransistorPmos: -3.84799e+07 muA
** NormalTransistorPmos: -3.84809e+07 muA
** NormalTransistorPmos: -3.84799e+07 muA
** NormalTransistorPmos: -3.84809e+07 muA
** NormalTransistorNmos: 7.69591e+07 muA
** DiodeTransistorNmos: 7.69601e+07 muA
** NormalTransistorNmos: 3.84791e+07 muA
** NormalTransistorNmos: 3.84791e+07 muA
** NormalTransistorNmos: 4.33211e+07 muA
** NormalTransistorNmos: 4.33201e+07 muA
** NormalTransistorPmos: -4.33219e+07 muA
** NormalTransistorPmos: -4.33209e+07 muA
** DiodeTransistorNmos: 4.33191e+07 muA
** DiodeTransistorNmos: 4.33181e+07 muA
** NormalTransistorPmos: -4.33199e+07 muA
** NormalTransistorPmos: -4.33209e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.51649e+07 muA


** Expected Voltages: 
** ibias: 1.24201  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceStageBiasComplementarySecondStage: 0.611001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 1.48201  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.622001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.86301  V
** innerStageBias: 0.865001  V
** innerTransconductance: 4.40001  V
** inner: 4.40001  V
** inner: 0.619001  V


.END