** Name: two_stage_single_output_op_amp_151_7

.MACRO two_stage_single_output_op_amp_151_7 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSimpleFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=5e-6
mMainBias3 ibias ibias sourceNmos sourceNmos nmos4 L=5e-6 W=12e-6
mMainBias4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=181e-6
mSimpleFirstStageLoad5 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSimpleFirstStageTransconductor6 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=63e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=5e-6 W=72e-6
mMainBias8 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=5e-6 W=146e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=5e-6 W=600e-6
mSimpleFirstStageLoad10 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=2e-6 W=5e-6
mSimpleFirstStageTransconductor11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=63e-6
mSimpleFirstStageLoad12 FirstStageYout1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=222e-6
mSecondStage1Transconductor13 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=448e-6
mSimpleFirstStageLoad14 outFirstStage inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=222e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 10.1001e-12
.EOM two_stage_single_output_op_amp_151_7

** Expected Performance Values: 
** Gain: 82 dB
** Power consumption: 4.63301 mW
** Area: 5767 (mu_m)^2
** Transit frequency: 6.25601 MHz
** Transit frequency with error factor: 6.23306 MHz
** Slew rate: 5.89631 V/mu_s
** Phase margin: 60.1606°
** CMRR: 91 dB
** VoutMax: 4.75 V
** VoutMin: 0.220001 V
** VcmMax: 5.21001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorNmos: 1.21697e+08 muA
** DiodeTransistorNmos: 1.16921e+08 muA
** NormalTransistorNmos: 1.16921e+08 muA
** NormalTransistorNmos: 1.16921e+08 muA
** DiodeTransistorNmos: 1.16921e+08 muA
** NormalTransistorPmos: -1.46918e+08 muA
** NormalTransistorPmos: -1.46918e+08 muA
** NormalTransistorNmos: 5.99951e+07 muA
** NormalTransistorNmos: 2.99981e+07 muA
** NormalTransistorNmos: 2.99981e+07 muA
** NormalTransistorNmos: 5.01139e+08 muA
** NormalTransistorPmos: -5.01138e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.21696e+08 muA


** Expected Voltages: 
** ibias: 0.626001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 4.24301  V
** out: 2.5  V
** outFirstStage: 4.18501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 1.15201  V
** innerTransistorStack1Load1: 1.15201  V
** out1: 2.30401  V
** sourceTransconductance: 1.94501  V


.END