** Name: two_stage_single_output_op_amp_68_9

.MACRO two_stage_single_output_op_amp_68_9 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=4e-6 W=6e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=13e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=278e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=33e-6
m5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=11e-6
m6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=167e-6
m7 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=4e-6 W=285e-6
m8 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=285e-6
m9 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=278e-6
m10 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=253e-6
m11 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=253e-6
m12 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=128e-6
m13 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=4e-6 W=128e-6
m14 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
m15 out outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=338e-6
m16 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=64e-6
m17 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=285e-6
m18 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=87e-6
m19 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourcePmos sourcePmos pmos4 L=4e-6 W=285e-6
m20 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=359e-6
m21 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=359e-6
m22 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=167e-6
m23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 13.6001e-12
.EOM two_stage_single_output_op_amp_68_9

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 11.6831 mW
** Area: 14999 (mu_m)^2
** Transit frequency: 5.14701 MHz
** Transit frequency with error factor: 5.14735 MHz
** Slew rate: 11.2036 V/mu_s
** Phase margin: 60.1606°
** CMRR: 139 dB
** VoutMax: 4.25 V
** VoutMin: 0.940001 V
** VcmMax: 3.07001 V
** VcmMin: -0.269999 V


** Expected Currents: 
** NormalTransistorPmos: -8.02089e+07 muA
** NormalTransistorPmos: -5.85549e+07 muA
** NormalTransistorNmos: 1.53968e+08 muA
** NormalTransistorNmos: 2.3095e+08 muA
** NormalTransistorNmos: 1.5397e+08 muA
** NormalTransistorNmos: 2.30952e+08 muA
** DiodeTransistorPmos: -1.53967e+08 muA
** NormalTransistorPmos: -1.53968e+08 muA
** NormalTransistorPmos: -1.53969e+08 muA
** DiodeTransistorPmos: -1.53968e+08 muA
** NormalTransistorPmos: -1.53965e+08 muA
** DiodeTransistorPmos: -1.53964e+08 muA
** NormalTransistorPmos: -7.69829e+07 muA
** NormalTransistorPmos: -7.69829e+07 muA
** NormalTransistorNmos: 1.71593e+09 muA
** DiodeTransistorNmos: 1.71593e+09 muA
** NormalTransistorPmos: -1.71592e+09 muA
** DiodeTransistorNmos: 8.02081e+07 muA
** NormalTransistorNmos: 8.02071e+07 muA
** DiodeTransistorNmos: 5.85541e+07 muA
** DiodeTransistorNmos: 5.85531e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.41801  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.77701  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.34801  V
** outSourceVoltageBiasXXnXX1: 0.674001  V
** outSourceVoltageBiasXXnXX2: 0.696001  V
** outSourceVoltageBiasXXpXX1: 4.21001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.08701  V
** innerTransistorStack2Load2: 4.08701  V
** out1: 3.34901  V
** sourceGCC1: 1.20201  V
** sourceGCC2: 1.20201  V
** sourceTransconductance: 3.40901  V
** inner: 0.672001  V
** inner: 4.20701  V


.END