** Name: two_stage_single_output_op_amp_31_8

.MACRO two_stage_single_output_op_amp_31_8 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=8e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
m3 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
m4 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=430e-6
m5 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=10e-6
m6 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=40e-6
m7 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=10e-6
m8 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=2e-6 W=41e-6
m9 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=600e-6
m10 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=155e-6
m11 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=79e-6
m12 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_31_8

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 3.24401 mW
** Area: 2615 (mu_m)^2
** Transit frequency: 4.44501 MHz
** Transit frequency with error factor: 4.44234 MHz
** Slew rate: 4.25176 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** negPSRR: 104 dB
** posPSRR: 98 dB
** VoutMax: 4.53001 V
** VoutMin: 0.740001 V
** VcmMax: 4.37001 V
** VcmMin: 1.27001 V


** Expected Currents: 
** NormalTransistorPmos: -1.96209e+07 muA
** NormalTransistorPmos: -1.96209e+07 muA
** DiodeTransistorPmos: -1.96209e+07 muA
** NormalTransistorNmos: 3.92391e+07 muA
** NormalTransistorNmos: 3.92401e+07 muA
** NormalTransistorNmos: 1.96201e+07 muA
** NormalTransistorNmos: 1.96201e+07 muA
** NormalTransistorNmos: 5.99612e+08 muA
** NormalTransistorNmos: 5.99611e+08 muA
** NormalTransistorPmos: -5.99611e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA


** Expected Voltages: 
** ibias: 1.13401  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.96901  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.578001  V
** innerTransistorStack2Load1: 4.13501  V
** out1: 3.40501  V
** sourceTransconductance: 1.94201  V
** innerStageBias: 0.547001  V


.END