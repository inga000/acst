** Name: symmetrical_op_amp79

.MACRO symmetrical_op_amp79 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=20e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias2 innerComplementarySecondStage innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=74e-6
mSymmetricalFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=600e-6
mMainBias4 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=8e-6 W=8e-6
mSecondStage1StageBias5 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mSymmetricalFirstStageLoad6 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=413e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=16e-6
mSymmetricalFirstStageLoad8 outFirstStage outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=413e-6
mSymmetricalFirstStageStageBias9 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=600e-6
mSecondStage1StageBias10 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=74e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=20e-6
mMainBias12 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=264e-6
mSymmetricalFirstStageTransconductor13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=99e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mSecondStage1StageBias15 out outVoltageBiasXXnXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=8e-6 W=259e-6
mSymmetricalFirstStageTransconductor16 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=99e-6
mSecondStage1Transconductor17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=555e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor18 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=555e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor19 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=142e-6
mSecondStage1Transconductor20 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=142e-6
mMainBias21 outVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=6e-6 W=49e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp79

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 4.32701 mW
** Area: 13893 (mu_m)^2
** Transit frequency: 10.6091 MHz
** Transit frequency with error factor: 10.6093 MHz
** Slew rate: 20.1485 V/mu_s
** Phase margin: 66.4632°
** CMRR: 143 dB
** negPSRR: 57 dB
** posPSRR: 44 dB
** VoutMax: 4.52001 V
** VoutMin: 0.450001 V
** VcmMax: 4.64001 V
** VcmMin: 1.41001 V


** Expected Currents: 
** NormalTransistorNmos: 5.50401e+06 muA
** NormalTransistorNmos: 1.31994e+08 muA
** NormalTransistorPmos: -1.69729e+07 muA
** DiodeTransistorPmos: -1.481e+08 muA
** DiodeTransistorPmos: -1.481e+08 muA
** NormalTransistorNmos: 2.962e+08 muA
** DiodeTransistorNmos: 2.96199e+08 muA
** NormalTransistorNmos: 1.48101e+08 muA
** NormalTransistorNmos: 1.48101e+08 muA
** NormalTransistorNmos: 2.0237e+08 muA
** NormalTransistorNmos: 2.02369e+08 muA
** NormalTransistorPmos: -2.02369e+08 muA
** NormalTransistorPmos: -2.02368e+08 muA
** DiodeTransistorNmos: 2.02368e+08 muA
** NormalTransistorPmos: -2.02367e+08 muA
** NormalTransistorPmos: -2.02368e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 1.69721e+07 muA
** DiodeTransistorPmos: -5.50499e+06 muA
** DiodeTransistorPmos: -1.31993e+08 muA


** Expected Voltages: 
** ibias: 1.11501  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 3.68601  V
** inSourceTransconductanceComplementarySecondStage: 4.23501  V
** innerComplementarySecondStage: 0.584001  V
** inputVoltageBiasXXpXX0: 4.09501  V
** out: 2.5  V
** outFirstStage: 4.23501  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outVoltageBiasXXnXX2: 0.855001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.79701  V
** innerStageBias: 0.179001  V
** innerTransconductance: 4.53101  V
** inner: 4.53101  V
** inner: 0.556001  V


.END