.suckt  two_stage_single_output_op_amp_182_2 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m3 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m5 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m6 outFirstStage FirstStageYinnerSourceLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m8 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m9 FirstStageYinnerTransistorStack1Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m11 FirstStageYinnerTransistorStack2Load2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m12 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m13 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m14 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c2 out sourceNmos 
m16 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m17 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m18 out ibias sourcePmos sourcePmos pmos
m19 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m20 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m21 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m23 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_182_2

