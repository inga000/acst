** Name: two_stage_single_output_op_amp_31_10

.MACRO two_stage_single_output_op_amp_31_10 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=4e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=11e-6
m3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m4 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=17e-6
m5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=9e-6 W=476e-6
m6 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=41e-6
m7 inputVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=4e-6 W=7e-6
m8 out ibias sourceNmos sourceNmos nmos4 L=4e-6 W=530e-6
m9 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=147e-6
m10 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=4e-6 W=45e-6
m11 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=5e-6 W=147e-6
m12 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=10e-6 W=83e-6
m13 out inputVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=600e-6
m14 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=124e-6
m15 outVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=49e-6
m16 FirstStageYout1 FirstStageYinnerTransistorStack2Load1 sourcePmos sourcePmos pmos4 L=9e-6 W=476e-6
m17 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=447e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 14.1001e-12
.EOM two_stage_single_output_op_amp_31_10

** Expected Performance Values: 
** Gain: 101 dB
** Power consumption: 7.97701 mW
** Area: 14931 (mu_m)^2
** Transit frequency: 8.38201 MHz
** Transit frequency with error factor: 8.37788 MHz
** Slew rate: 7.89989 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** negPSRR: 108 dB
** posPSRR: 101 dB
** VoutMax: 4.25 V
** VoutMin: 0.340001 V
** VcmMax: 4.44001 V
** VcmMin: 1.70001 V


** Expected Currents: 
** NormalTransistorNmos: 1.72201e+07 muA
** NormalTransistorNmos: 1.01534e+08 muA
** NormalTransistorPmos: -5.04859e+07 muA
** NormalTransistorPmos: -5.59969e+07 muA
** NormalTransistorPmos: -5.59969e+07 muA
** DiodeTransistorPmos: -5.59969e+07 muA
** NormalTransistorNmos: 1.11992e+08 muA
** NormalTransistorNmos: 1.11991e+08 muA
** NormalTransistorNmos: 5.59961e+07 muA
** NormalTransistorNmos: 5.59961e+07 muA
** NormalTransistorNmos: 1.30407e+09 muA
** NormalTransistorPmos: -1.30406e+09 muA
** NormalTransistorPmos: -1.30406e+09 muA
** DiodeTransistorNmos: 5.04851e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.72209e+07 muA
** DiodeTransistorPmos: -1.01533e+08 muA


** Expected Voltages: 
** ibias: 0.747001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 3.95801  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 4.03301  V
** outVoltageBiasXXnXX1: 1.14501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.342001  V
** innerTransistorStack2Load1: 4.19201  V
** out1: 3.46901  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.59701  V


.END