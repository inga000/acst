** Name: two_stage_single_output_op_amp_167_3

.MACRO two_stage_single_output_op_amp_167_3 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=60e-6
m2 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=24e-6
m3 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m4 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=544e-6
m5 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=4e-6 W=478e-6
m6 outFirstStage outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=324e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=496e-6
m8 FirstStageYout1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=324e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=478e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=77e-6
m11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=598e-6
m12 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=73e-6
m13 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
m14 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=4e-6 W=544e-6
m15 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=77e-6
m16 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=45e-6
m17 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=311e-6
Capacitor1 outFirstStage out 6.5e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_167_3

** Expected Performance Values: 
** Gain: 80 dB
** Power consumption: 6.06601 mW
** Area: 14764 (mu_m)^2
** Transit frequency: 4.39701 MHz
** Transit frequency with error factor: 4.35424 MHz
** Slew rate: 5.58641 V/mu_s
** Phase margin: 60.1606°
** CMRR: 96 dB
** VoutMax: 4.03001 V
** VoutMin: 0.150001 V
** VcmMax: 3.22001 V
** VcmMin: -0.289999 V


** Expected Currents: 
** NormalTransistorPmos: -7.33199e+07 muA
** DiodeTransistorPmos: -3.8357e+08 muA
** DiodeTransistorPmos: -3.83571e+08 muA
** NormalTransistorPmos: -3.8357e+08 muA
** NormalTransistorPmos: -3.83571e+08 muA
** NormalTransistorNmos: 4.02328e+08 muA
** NormalTransistorNmos: 4.02328e+08 muA
** NormalTransistorPmos: -3.75139e+07 muA
** NormalTransistorPmos: -3.75129e+07 muA
** NormalTransistorPmos: -1.87569e+07 muA
** NormalTransistorPmos: -1.87569e+07 muA
** NormalTransistorNmos: 3.15317e+08 muA
** NormalTransistorPmos: -3.15316e+08 muA
** NormalTransistorPmos: -3.15315e+08 muA
** DiodeTransistorNmos: 7.33191e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.48201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.675001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 4.03701  V
** innerStageBias: 4.26101  V
** innerTransistorStack2Load1: 4.03401  V
** out1: 3.04801  V
** sourceTransconductance: 3.26601  V
** innerStageBias: 4.21701  V


.END