** Name: two_stage_single_output_op_amp_55_1

.MACRO two_stage_single_output_op_amp_55_1 ibias in1 in2 out sourceNmos sourcePmos
m1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=57e-6
m2 ibias ibias sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
m3 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=57e-6
m4 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
m5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=6e-6
m6 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=57e-6
m7 outVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=88e-6
m8 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=2e-6 W=24e-6
m9 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=57e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=36e-6
m11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=2e-6 W=72e-6
m12 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=2e-6 W=36e-6
m13 out outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=442e-6
m14 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=316e-6
m15 FirstStageYsourceGCC1 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
m16 FirstStageYsourceGCC2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
m17 out outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=587e-6
m18 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=316e-6
Capacitor1 outFirstStage out 17.3001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_55_1

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 9.13501 mW
** Area: 6626 (mu_m)^2
** Transit frequency: 4.74901 MHz
** Transit frequency with error factor: 4.74899 MHz
** Slew rate: 3.69268 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.63001 V
** VoutMin: 0.560001 V
** VcmMax: 5.03001 V
** VcmMin: 0.75 V


** Expected Currents: 
** NormalTransistorNmos: 3.00031e+07 muA
** NormalTransistorNmos: 1.07834e+08 muA
** NormalTransistorPmos: -6.41689e+07 muA
** NormalTransistorPmos: -1.08283e+08 muA
** NormalTransistorPmos: -6.41689e+07 muA
** NormalTransistorPmos: -1.08283e+08 muA
** DiodeTransistorNmos: 6.41681e+07 muA
** NormalTransistorNmos: 6.41671e+07 muA
** NormalTransistorNmos: 6.41681e+07 muA
** DiodeTransistorNmos: 6.41671e+07 muA
** NormalTransistorNmos: 8.82271e+07 muA
** NormalTransistorNmos: 4.41141e+07 muA
** NormalTransistorNmos: 4.41141e+07 muA
** NormalTransistorNmos: 1.46256e+09 muA
** NormalTransistorPmos: -1.46255e+09 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -3.00039e+07 muA
** DiodeTransistorPmos: -1.07833e+08 muA


** Expected Voltages: 
** ibias: 0.576001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.967001  V
** outVoltageBiasXXpXX1: 3.68601  V
** outVoltageBiasXXpXX2: 4.06101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.604001  V
** innerTransistorStack1Load2: 0.604001  V
** out1: 1.17201  V
** sourceGCC1: 4.40001  V
** sourceGCC2: 4.40001  V
** sourceTransconductance: 1.92401  V


.END