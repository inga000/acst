.suckt  two_stage_single_output_op_amp_156_3 ibias in1 in2 out sourceNmos sourcePmos
cCompensationCapacitor1 outFirstStage out 
mMainBias1 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
mMainBias2 outInputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad3 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad4 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos
mSimpleFirstStageLoad5 FirstStageYout1 ibias sourceNmos sourceNmos nmos
mSimpleFirstStageLoad6 outFirstStage ibias sourceNmos sourceNmos nmos
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
mSimpleFirstStageStageBias8 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
cLoadCapacitor2 out sourceNmos 
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos
mSecondStage1StageBias12 out outInputVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
mSecondStage1StageBias13 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
mMainBias14 ibias ibias sourceNmos sourceNmos nmos
mMainBias15 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
mMainBias17 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
mMainBias18 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_156_3

