** Name: two_stage_single_output_op_amp_1_5

.MACRO two_stage_single_output_op_amp_1_5 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=143e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=14e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=21e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=67e-6
mSecondStage1Transconductor6 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=188e-6
mSimpleFirstStageLoad7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=143e-6
mMainBias8 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=1e-6 W=13e-6
mSimpleFirstStageTransconductor9 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=25e-6
mSimpleFirstStageStageBias10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=60e-6
mMainBias11 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=21e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=67e-6
mSimpleFirstStageTransconductor13 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=25e-6
mMainBias14 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=41e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_1_5

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 1.40301 mW
** Area: 4380 (mu_m)^2
** Transit frequency: 2.87901 MHz
** Transit frequency with error factor: 2.8632 MHz
** Slew rate: 4.88521 V/mu_s
** Phase margin: 67.6091°
** CMRR: 87 dB
** negPSRR: 89 dB
** posPSRR: 199 dB
** VoutMax: 3.16001 V
** VoutMin: 0.150001 V
** VcmMax: 3.46001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 3.83301e+07 muA
** NormalTransistorPmos: -4.15689e+07 muA
** DiodeTransistorNmos: 3.04151e+07 muA
** NormalTransistorNmos: 3.04151e+07 muA
** NormalTransistorPmos: -6.08319e+07 muA
** NormalTransistorPmos: -3.04159e+07 muA
** NormalTransistorPmos: -3.04159e+07 muA
** NormalTransistorNmos: 1.19966e+08 muA
** NormalTransistorPmos: -1.19965e+08 muA
** DiodeTransistorPmos: -1.19966e+08 muA
** DiodeTransistorNmos: 4.15681e+07 muA
** DiodeTransistorPmos: -3.83309e+07 muA
** NormalTransistorPmos: -3.83319e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.19901  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 2.60001  V
** outSourceVoltageBiasXXpXX1: 3.80001  V
** outVoltageBiasXXnXX0: 0.592001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceTransconductance: 3.79901  V
** inner: 3.80001  V


.END