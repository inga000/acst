** Name: symmetrical_op_amp51

.MACRO symmetrical_op_amp51 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=8e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=8e-6 W=63e-6
mMainBias3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=6e-6
mSymmetricalFirstStageLoad4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=63e-6
mMainBias5 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=4e-6 W=40e-6
mMainBias6 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=8e-6
mSymmetricalFirstStageStageBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=157e-6
mSecondStage1Transconductor8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=8e-6 W=137e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=8e-6 W=137e-6
mMainBias10 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=14e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor11 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=32e-6
mSecondStage1Transconductor12 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=32e-6
mSymmetricalFirstStageStageBias13 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=157e-6
mSecondStage1StageBias14 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=260e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias15 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=260e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=40e-6
mMainBias17 inOutputTransconductanceComplementarySecondStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=102e-6
mSymmetricalFirstStageTransconductor18 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=46e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias19 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=4e-6 W=35e-6
mMainBias20 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=34e-6
mSecondStage1StageBias21 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=4e-6 W=342e-6
mSymmetricalFirstStageTransconductor22 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=3e-6 W=46e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp51

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 0.996001 mW
** Area: 9768 (mu_m)^2
** Transit frequency: 2.54501 MHz
** Transit frequency with error factor: 2.54537 MHz
** Slew rate: 4.22938 V/mu_s
** Phase margin: 62.4525°
** CMRR: 146 dB
** negPSRR: 45 dB
** posPSRR: 50 dB
** VoutMax: 4.64001 V
** VoutMin: 0.480001 V
** VcmMax: 3.13001 V
** VcmMin: 0.0100001 V


** Expected Currents: 
** NormalTransistorNmos: 2.03051e+07 muA
** NormalTransistorPmos: -8.61699e+06 muA
** NormalTransistorPmos: -2.55339e+07 muA
** DiodeTransistorNmos: 1.98961e+07 muA
** DiodeTransistorNmos: 1.98961e+07 muA
** NormalTransistorPmos: -3.97949e+07 muA
** DiodeTransistorPmos: -3.97939e+07 muA
** NormalTransistorPmos: -1.98969e+07 muA
** NormalTransistorPmos: -1.98969e+07 muA
** NormalTransistorNmos: 4.24611e+07 muA
** NormalTransistorNmos: 4.24621e+07 muA
** NormalTransistorPmos: -4.24619e+07 muA
** NormalTransistorPmos: -4.24629e+07 muA
** NormalTransistorPmos: -4.24639e+07 muA
** NormalTransistorPmos: -4.24649e+07 muA
** NormalTransistorNmos: 4.24631e+07 muA
** NormalTransistorNmos: 4.24621e+07 muA
** DiodeTransistorNmos: 8.61601e+06 muA
** DiodeTransistorNmos: 2.55331e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -2.03059e+07 muA


** Expected Voltages: 
** ibias: 3.39601  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 3.68601  V
** inOutputTransconductanceComplementarySecondStage: 0.883001  V
** inSourceTransconductanceComplementarySecondStage: 0.577001  V
** innerComplementarySecondStage: 4.24401  V
** inputVoltageBiasXXnXX0: 0.725001  V
** out: 2.5  V
** outFirstStage: 0.577001  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.33301  V
** innerStageBias: 4.41601  V
** innerTransconductance: 0.172001  V
** inner: 4.76901  V
** inner: 0.172001  V
** inner: 4.19601  V


.END