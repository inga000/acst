** Name: two_stage_single_output_op_amp_4_2

.MACRO two_stage_single_output_op_amp_4_2 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=27e-6
m2 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 nmos4 L=8e-6 W=128e-6
m3 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=67e-6
m4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=11e-6
m5 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=533e-6
m6 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=8e-6 W=128e-6
m7 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=8e-6 W=67e-6
m8 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=281e-6
m9 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=1e-6 W=283e-6
m10 out ibias sourcePmos sourcePmos pmos4 L=1e-6 W=589e-6
m11 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=29e-6
m12 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=29e-6
m13 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=107e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_4_2

** Expected Performance Values: 
** Gain: 85 dB
** Power consumption: 4.61301 mW
** Area: 9111 (mu_m)^2
** Transit frequency: 5.34201 MHz
** Transit frequency with error factor: 5.32504 MHz
** Slew rate: 20.709 V/mu_s
** Phase margin: 60.1606°
** CMRR: 92 dB
** negPSRR: 93 dB
** posPSRR: 109 dB
** VoutMax: 4.77001 V
** VoutMin: 0.670001 V
** VcmMax: 3.60001 V
** VcmMin: 0.700001 V


** Expected Currents: 
** NormalTransistorPmos: -2.6091e+08 muA
** DiodeTransistorNmos: 4.93231e+07 muA
** DiodeTransistorNmos: 4.93221e+07 muA
** NormalTransistorNmos: 4.93231e+07 muA
** NormalTransistorNmos: 4.93221e+07 muA
** NormalTransistorPmos: -9.86479e+07 muA
** NormalTransistorPmos: -4.93239e+07 muA
** NormalTransistorPmos: -4.93239e+07 muA
** NormalTransistorNmos: 5.43027e+08 muA
** NormalTransistorNmos: 5.43026e+08 muA
** NormalTransistorPmos: -5.43026e+08 muA
** DiodeTransistorNmos: 2.60911e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.21001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.07801  V
** out: 2.5  V
** outFirstStage: 0.858001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 1.26301  V
** innerSourceLoad1: 0.668001  V
** innerTransistorStack2Load1: 0.667001  V
** sourceTransconductance: 3.67801  V
** innerTransconductance: 0.453001  V


.END