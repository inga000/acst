** Name: symmetrical_op_amp149

.MACRO symmetrical_op_amp149 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=14e-6
m2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=21e-6
m3 innerComplementarySecondStage innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=174e-6
m4 ibias ibias VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=13e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=43e-6
m6 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=8e-6 W=49e-6
m7 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=7e-6 W=19e-6
m8 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=7e-6 W=61e-6
m9 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=7e-6 W=19e-6
m10 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=7e-6 W=61e-6
m11 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=2e-6 W=33e-6
m12 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=51e-6
m13 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=51e-6
m14 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=7e-6 W=113e-6
m15 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=7e-6 W=113e-6
m16 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=239e-6
m17 out outVoltageBiasXXpXX2 SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=8e-6 W=583e-6
m18 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=239e-6
m19 out2FirstStage outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=69e-6
m20 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=52e-6
m21 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=43e-6
m22 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=7e-6 W=174e-6
m23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=13e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp149

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 1.41601 mW
** Area: 14926 (mu_m)^2
** Transit frequency: 3.54501 MHz
** Transit frequency with error factor: 3.54474 MHz
** Slew rate: 3.66015 V/mu_s
** Phase margin: 60.1606°
** CMRR: 149 dB
** negPSRR: 46 dB
** posPSRR: 49 dB
** VoutMax: 4.54001 V
** VoutMin: 0.560001 V
** VcmMax: 3.12001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorNmos: 6.21881e+07 muA
** NormalTransistorPmos: -4.03509e+07 muA
** NormalTransistorPmos: -5.34559e+07 muA
** NormalTransistorNmos: 1.67721e+07 muA
** NormalTransistorNmos: 1.67711e+07 muA
** NormalTransistorNmos: 1.67721e+07 muA
** NormalTransistorNmos: 1.67711e+07 muA
** NormalTransistorPmos: -3.35449e+07 muA
** DiodeTransistorPmos: -3.35439e+07 muA
** NormalTransistorPmos: -1.67729e+07 muA
** NormalTransistorPmos: -1.67729e+07 muA
** NormalTransistorNmos: 3.68341e+07 muA
** NormalTransistorNmos: 3.68351e+07 muA
** NormalTransistorPmos: -3.68349e+07 muA
** NormalTransistorPmos: -3.68359e+07 muA
** DiodeTransistorPmos: -3.68349e+07 muA
** NormalTransistorNmos: 3.68341e+07 muA
** NormalTransistorNmos: 3.68351e+07 muA
** DiodeTransistorNmos: 4.03501e+07 muA
** DiodeTransistorNmos: 5.34551e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** NormalTransistorPmos: -1e+07 muA
** DiodeTransistorPmos: -6.21889e+07 muA


** Expected Voltages: 
** ibias: 3.28201  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.570001  V
** innerComplementarySecondStage: 4.14701  V
** out: 2.5  V
** out1FirstStage: 0.570001  V
** out2FirstStage: 0.969001  V
** outSourceVoltageBiasXXpXX1: 4.14201  V
** outVoltageBiasXXnXX0: 0.617001  V
** outVoltageBiasXXpXX2: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.413001  V
** innerTransistorStack2Load1: 0.413001  V
** sourceTransconductance: 3.22901  V
** innerStageBias: 4.41801  V
** innerTransconductance: 0.165001  V
** inner: 0.165001  V
** inner: 4.13801  V


.END