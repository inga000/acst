** Name: two_stage_single_output_op_amp_43_8

.MACRO two_stage_single_output_op_amp_43_8 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=9e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=8e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=114e-6
m4 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=88e-6
m5 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=2e-6 W=161e-6
m6 outFirstStage inputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=44e-6
m7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=44e-6
m8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=58e-6
m9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=58e-6
m10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=209e-6
m11 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=103e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=475e-6
m13 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=1e-6 W=88e-6
m14 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=326e-6
m15 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=7e-6 W=326e-6
m16 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=7e-6 W=549e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10.4001e-12
.EOM two_stage_single_output_op_amp_43_8

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 2.01101 mW
** Area: 11759 (mu_m)^2
** Transit frequency: 4.35601 MHz
** Transit frequency with error factor: 4.35037 MHz
** Slew rate: 4.01657 V/mu_s
** Phase margin: 60.1606°
** CMRR: 105 dB
** VoutMax: 4.83001 V
** VoutMin: 0.760001 V
** VcmMax: 4.08001 V
** VcmMin: -0.399999 V


** Expected Currents: 
** NormalTransistorPmos: -9.01699e+06 muA
** NormalTransistorNmos: 4.19021e+07 muA
** NormalTransistorNmos: 6.63891e+07 muA
** NormalTransistorNmos: 4.19021e+07 muA
** NormalTransistorNmos: 6.63891e+07 muA
** DiodeTransistorPmos: -4.19029e+07 muA
** NormalTransistorPmos: -4.19029e+07 muA
** NormalTransistorPmos: -4.89759e+07 muA
** NormalTransistorPmos: -2.44879e+07 muA
** NormalTransistorPmos: -2.44879e+07 muA
** NormalTransistorNmos: 2.40325e+08 muA
** NormalTransistorNmos: 2.40324e+08 muA
** NormalTransistorPmos: -2.40324e+08 muA
** DiodeTransistorNmos: 9.01601e+06 muA
** DiodeTransistorNmos: 9.01701e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.12801  V
** out: 2.5  V
** outFirstStage: 4.26701  V
** outSourceVoltageBiasXXnXX1: 0.569001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 4.27201  V
** sourceGCC1: 0.573001  V
** sourceGCC2: 0.573001  V
** sourceTransconductance: 3.23501  V
** innerStageBias: 0.535001  V


.END