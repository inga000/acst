.suckt  complementary_op_amp1 ibias in1 in2 out sourceNmos sourcePmos
m_Complementary_MainBias_1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_2 FirstStageYinnerOutputLoadPmos FirstStageYinnerOutputLoadPmos FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos pmos
m_Complementary_FirstStage_Load_3 FirstStageYinnerSourceLoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_4 out FirstStageYinnerOutputLoadPmos FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerTransistorStack2LoadPmos pmos
m_Complementary_FirstStage_Load_5 FirstStageYinnerTransistorStack2LoadPmos FirstStageYinnerSourceLoadPmos sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Load_6 FirstStageYinnerOutputLoadPmos FirstStageYinnerOutputLoadPmos FirstStageYinnerSourceLoadNmos FirstStageYinnerSourceLoadNmos nmos
m_Complementary_FirstStage_Load_7 FirstStageYinnerSourceLoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_Load_8 out FirstStageYinnerOutputLoadPmos FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerTransistorStack2LoadNmos nmos
m_Complementary_FirstStage_Load_9 FirstStageYinnerTransistorStack2LoadNmos FirstStageYinnerSourceLoadNmos sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_10 FirstStageYsourceTransconductanceNmos outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_FirstStage_StageBias_11 FirstStageYsourceTransconductancePmos ibias sourcePmos sourcePmos pmos
m_Complementary_FirstStage_Transconductor_12 FirstStageYinnerSourceLoadPmos in1 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_13 FirstStageYinnerTransistorStack2LoadPmos in2 FirstStageYsourceTransconductanceNmos FirstStageYsourceTransconductanceNmos nmos
m_Complementary_FirstStage_Transconductor_14 FirstStageYinnerSourceLoadNmos in1 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
m_Complementary_FirstStage_Transconductor_15 FirstStageYinnerTransistorStack2LoadNmos in2 FirstStageYsourceTransconductancePmos FirstStageYsourceTransconductancePmos pmos
c_Complementary_Load_Capacitor_1 out sourceNmos 
m_Complementary_MainBias_16 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_Complementary_MainBias_17 ibias ibias sourcePmos sourcePmos pmos
.end complementary_op_amp1

