** Name: one_stage_single_output_op_amp79

.MACRO one_stage_single_output_op_amp79 ibias in1 in2 out sourceNmos sourcePmos
m1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=51e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=5e-6 W=7e-6
m3 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=23e-6
m4 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m5 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=5e-6 W=128e-6
m6 FirstStageYinnerStageBias inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=210e-6
m7 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=135e-6
m8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=5e-6 W=135e-6
m9 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=5e-6 W=128e-6
m10 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=15e-6
m11 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=15e-6
m12 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=5e-6 W=156e-6
m13 out ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=124e-6
m14 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
m15 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=37e-6
m16 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=124e-6
m17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=107e-6
m18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=107e-6
Capacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp79

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 1.45801 mW
** Area: 5851 (mu_m)^2
** Transit frequency: 3.40101 MHz
** Transit frequency with error factor: 3.40066 MHz
** Slew rate: 3.60577 V/mu_s
** Phase margin: 88.8085°
** CMRR: 145 dB
** VoutMax: 4.02001 V
** VoutMin: 0.360001 V
** VcmMax: 5.17001 V
** VcmMin: 1.31001 V


** Expected Currents: 
** NormalTransistorPmos: -3.74069e+07 muA
** NormalTransistorPmos: -1.72349e+07 muA
** NormalTransistorPmos: -7.23229e+07 muA
** NormalTransistorPmos: -1.08482e+08 muA
** NormalTransistorPmos: -7.23249e+07 muA
** NormalTransistorPmos: -1.08484e+08 muA
** NormalTransistorNmos: 7.23221e+07 muA
** NormalTransistorNmos: 7.23231e+07 muA
** NormalTransistorNmos: 7.23241e+07 muA
** NormalTransistorNmos: 7.23231e+07 muA
** NormalTransistorNmos: 7.23211e+07 muA
** NormalTransistorNmos: 7.23201e+07 muA
** NormalTransistorNmos: 3.61611e+07 muA
** NormalTransistorNmos: 3.61611e+07 muA
** DiodeTransistorNmos: 3.74061e+07 muA
** DiodeTransistorNmos: 1.72351e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.47901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 0.573001  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX1: 0.964001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.393001  V
** innerTransistorStack1Load2: 0.376001  V
** innerTransistorStack2Load2: 0.377001  V
** out1: 0.582001  V
** sourceGCC1: 4.22301  V
** sourceGCC2: 4.22301  V
** sourceTransconductance: 1.92601  V


.END