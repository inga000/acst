.suckt  two_stage_fully_differential_op_amp_44_6 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c1 out1FirstStage out1 
c2 out2FirstStage out2 
m1 outInputVoltageBiasXXpXX1 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m2 outInputVoltageBiasXXpXX2 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m3 outInputVoltageBiasXXpXX3 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m4 outVoltageBiasXXpXX4 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m5 inputVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX5 sourcePmos sourcePmos pmos
m6 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX5 sourcePmos sourcePmos pmos
m7 FeedbackStageYout1 FeedbackStageYout1 sourceNmos sourceNmos nmos
m8 outFeedback outFeedback sourceNmos sourceNmos nmos
m9 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 pmos
m10 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXpXX5 sourcePmos sourcePmos pmos
m11 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 pmos
m12 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXpXX5 sourcePmos sourcePmos pmos
m13 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m14 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 pmos
m15 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m16 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 pmos
m17 out1FirstStage outVoltageBiasXXpXX4 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos
m18 out2FirstStage outVoltageBiasXXpXX4 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos
m19 out1FirstStage outFeedback sourceNmos sourceNmos nmos
m20 out2FirstStage outFeedback sourceNmos sourceNmos nmos
m21 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m22 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m23 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos
m24 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos
c3 out1 sourceNmos 
c4 out2 sourceNmos 
m25 out1 outVoltageBiasXXnXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance nmos
m26 SecondStage1YinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m27 out1 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos
m28 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m29 out2 outVoltageBiasXXnXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance nmos
m30 SecondStage2YinnerTransconductance out2FirstStage sourceNmos sourceNmos nmos
m31 out2 outInputVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 pmos
m32 outSourceVoltageBiasXXpXX3 outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m33 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos
m34 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m35 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m36 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m37 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos
m38 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m39 outInputVoltageBiasXXpXX3 outInputVoltageBiasXXpXX3 VoltageBiasXXpXX3Yinner VoltageBiasXXpXX3Yinner pmos
m40 VoltageBiasXXpXX3Yinner outSourceVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m41 outVoltageBiasXXpXX4 outVoltageBiasXXpXX4 sourceTransconductance sourceTransconductance pmos
m42 ibias ibias outSourceVoltageBiasXXpXX5 outSourceVoltageBiasXXpXX5 pmos
m43 outSourceVoltageBiasXXpXX5 outSourceVoltageBiasXXpXX5 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_44_6

