** Name: symmetrical_op_amp193

.MACRO symmetrical_op_amp193 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=3e-6 W=8e-6
mMainBias2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=17e-6
mSymmetricalFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=273e-6
mMainBias4 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=12e-6
mMainBias5 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=16e-6
mSymmetricalFirstStageStageBias6 FirstStageYsourceTransconductance ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=3e-6 W=273e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=104e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias8 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=104e-6
mMainBias9 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mSymmetricalFirstStageTransconductor10 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=103e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias11 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=1e-6 W=53e-6
mSecondStage1StageBias12 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=53e-6
mSymmetricalFirstStageTransconductor13 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=9e-6 W=103e-6
mMainBias14 out2FirstStage outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=98e-6
mMainBias15 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=18e-6
mSymmetricalFirstStageLoad16 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=104e-6
mSymmetricalFirstStageLoad17 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=104e-6
mSecondStage1Transconductor18 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=4e-6 W=129e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor19 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=4e-6 W=129e-6
mMainBias20 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=4e-6 W=143e-6
mSymmetricalFirstStageLoad21 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=415e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor22 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=1e-6 W=516e-6
mSecondStage1Transconductor23 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=1e-6 W=516e-6
mSymmetricalFirstStageLoad24 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=1e-6 W=415e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp193

** Expected Performance Values: 
** Gain: 92 dB
** Power consumption: 5.52301 mW
** Area: 8593 (mu_m)^2
** Transit frequency: 7.92001 MHz
** Transit frequency with error factor: 7.92021 MHz
** Slew rate: 20.8301 V/mu_s
** Phase margin: 81.933°
** CMRR: 134 dB
** negPSRR: 117 dB
** posPSRR: 56 dB
** VoutMax: 4.25 V
** VoutMin: 0.370001 V
** VcmMax: 4.81001 V
** VcmMin: 1.65001 V


** Expected Currents: 
** NormalTransistorNmos: 2.22391e+07 muA
** NormalTransistorNmos: 1.2184e+08 muA
** NormalTransistorPmos: -1.95056e+08 muA
** NormalTransistorPmos: -1.68172e+08 muA
** NormalTransistorPmos: -1.68173e+08 muA
** NormalTransistorPmos: -1.68172e+08 muA
** NormalTransistorPmos: -1.68173e+08 muA
** NormalTransistorNmos: 3.36346e+08 muA
** DiodeTransistorNmos: 3.36347e+08 muA
** NormalTransistorNmos: 1.68173e+08 muA
** NormalTransistorNmos: 1.68173e+08 muA
** NormalTransistorNmos: 2.09566e+08 muA
** NormalTransistorNmos: 2.09565e+08 muA
** NormalTransistorPmos: -2.09565e+08 muA
** NormalTransistorPmos: -2.09565e+08 muA
** NormalTransistorNmos: 2.09566e+08 muA
** NormalTransistorNmos: 2.09565e+08 muA
** NormalTransistorPmos: -2.09565e+08 muA
** NormalTransistorPmos: -2.09565e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 1.95057e+08 muA
** DiodeTransistorPmos: -2.22399e+07 muA
** DiodeTransistorPmos: -1.21839e+08 muA


** Expected Voltages: 
** ibias: 1.22801  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.775001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.559001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outSourceVoltageBiasXXnXX1: 0.615001  V
** outVoltageBiasXXpXX0: 3.88101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.67701  V
** innerStageBias: 0.154001  V
** innerTransconductance: 4.40001  V
** inner: 0.154001  V
** inner: 4.40001  V
** inner: 0.612001  V


.END