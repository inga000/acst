** Name: two_stage_single_output_op_amp_46_7

.MACRO two_stage_single_output_op_amp_46_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=22e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=19e-6
m4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=164e-6
m5 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=325e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=564e-6
m7 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=7e-6 W=530e-6
m8 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=7e-6 W=530e-6
m9 FirstStageYsourceGCC1 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=88e-6
m10 FirstStageYsourceGCC2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=88e-6
m11 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=145e-6
m12 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=325e-6
m13 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=102e-6
m14 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=106e-6
m15 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=1e-6 W=164e-6
m16 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=84e-6
m17 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=84e-6
m18 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=3e-6 W=308e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 18.8001e-12
.EOM two_stage_single_output_op_amp_46_7

** Expected Performance Values: 
** Gain: 114 dB
** Power consumption: 10.2761 mW
** Area: 14686 (mu_m)^2
** Transit frequency: 2.94401 MHz
** Transit frequency with error factor: 2.94377 MHz
** Slew rate: 7.58965 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 4.25 V
** VoutMin: 0.390001 V
** VcmMax: 3.67001 V
** VcmMin: -0.169999 V


** Expected Currents: 
** NormalTransistorPmos: -5.36569e+07 muA
** NormalTransistorPmos: -5.63799e+07 muA
** NormalTransistorNmos: 1.44211e+08 muA
** NormalTransistorNmos: 2.26495e+08 muA
** NormalTransistorNmos: 1.44209e+08 muA
** NormalTransistorNmos: 2.26493e+08 muA
** DiodeTransistorPmos: -1.4421e+08 muA
** DiodeTransistorPmos: -1.44209e+08 muA
** NormalTransistorPmos: -1.44208e+08 muA
** NormalTransistorPmos: -1.44209e+08 muA
** NormalTransistorPmos: -1.64569e+08 muA
** NormalTransistorPmos: -8.22849e+07 muA
** NormalTransistorPmos: -8.22849e+07 muA
** NormalTransistorNmos: 1.47225e+09 muA
** NormalTransistorPmos: -1.47224e+09 muA
** DiodeTransistorNmos: 5.36561e+07 muA
** DiodeTransistorNmos: 5.63791e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outVoltageBiasXXnXX1: 1.14601  V
** outVoltageBiasXXnXX2: 0.796001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.21401  V
** innerTransistorStack2Load2: 4.21301  V
** out1: 3.49201  V
** sourceGCC1: 0.591001  V
** sourceGCC2: 0.591001  V
** sourceTransconductance: 3.53001  V


.END