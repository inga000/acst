** Name: two_stage_single_output_op_amp_52_9

.MACRO two_stage_single_output_op_amp_52_9 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=28e-6
mMainBias2 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=9e-6 W=51e-6
mMainBias3 inputVoltageBiasXXnXX3 inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias4 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias5 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=525e-6
mMainBias6 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=7e-6 W=114e-6
mMainBias7 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=30e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=7e-6 W=28e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=5e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=5e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance inputVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=3e-6 W=19e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mSecondStage1StageBias13 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=525e-6
mFoldedCascodeFirstStageLoad14 outFirstStage inputVoltageBiasXXnXX2 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=9e-6 W=81e-6
mFoldedCascodeFirstStageLoad15 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=7e-6 W=172e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=90e-6
mFoldedCascodeFirstStageLoad17 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=90e-6
mMainBias18 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=522e-6
mMainBias19 inputVoltageBiasXXnXX3 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=13e-6
mSecondStage1Transconductor20 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=263e-6
mFoldedCascodeFirstStageLoad21 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=7e-6 W=172e-6
mMainBias22 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=7e-6 W=76e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_52_9

** Expected Performance Values: 
** Gain: 119 dB
** Power consumption: 14.7841 mW
** Area: 13015 (mu_m)^2
** Transit frequency: 2.64301 MHz
** Transit frequency with error factor: 2.64252 MHz
** Slew rate: 4.46284 V/mu_s
** Phase margin: 61.3065°
** CMRR: 137 dB
** VoutMax: 4.25 V
** VoutMin: 1.09001 V
** VcmMax: 5.04001 V
** VcmMin: 0.870001 V


** Expected Currents: 
** NormalTransistorPmos: -2.54449e+07 muA
** NormalTransistorPmos: -1.75566e+08 muA
** NormalTransistorPmos: -4.33599e+06 muA
** NormalTransistorPmos: -2.03869e+07 muA
** NormalTransistorPmos: -3.05799e+07 muA
** NormalTransistorPmos: -2.03869e+07 muA
** NormalTransistorPmos: -3.05799e+07 muA
** DiodeTransistorNmos: 2.03861e+07 muA
** NormalTransistorNmos: 2.03861e+07 muA
** NormalTransistorNmos: 2.03861e+07 muA
** NormalTransistorNmos: 2.03871e+07 muA
** NormalTransistorNmos: 1.01941e+07 muA
** NormalTransistorNmos: 1.01941e+07 muA
** NormalTransistorNmos: 2.67035e+09 muA
** DiodeTransistorNmos: 2.67035e+09 muA
** NormalTransistorPmos: -2.67034e+09 muA
** DiodeTransistorNmos: 2.54441e+07 muA
** NormalTransistorNmos: 2.54431e+07 muA
** DiodeTransistorNmos: 1.75567e+08 muA
** DiodeTransistorNmos: 4.33501e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.01301  V
** inputVoltageBiasXXnXX3: 0.600001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.5  V
** outSourceVoltageBiasXXnXX1: 0.75  V
** outSourceVoltageBiasXXpXX1: 4.07301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.445001  V
** out1: 0.650001  V
** sourceGCC1: 4.10201  V
** sourceGCC2: 4.10201  V
** sourceTransconductance: 1.82501  V
** inner: 0.747001  V


.END