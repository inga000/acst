** Name: symmetrical_op_amp97

.MACRO symmetrical_op_amp97 ibias in1 in2 out sourceNmos sourcePmos
m1 out2FirstStage out2FirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
m2 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=89e-6
m3 inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
m4 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=2e-6 W=23e-6
m5 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=2e-6 W=18e-6
m6 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=2e-6 W=18e-6
m7 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos4 L=2e-6 W=23e-6
m8 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
m9 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
m10 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
m11 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=1e-6 W=20e-6
m12 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=90e-6
m13 innerComplementarySecondStage inStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=44e-6
m14 out innerComplementarySecondStage inStageBiasComplementarySecondStage inStageBiasComplementarySecondStage pmos4 L=1e-6 W=48e-6
m15 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=90e-6
m16 out2FirstStage ibias sourcePmos sourcePmos pmos4 L=6e-6 W=260e-6
m17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=600e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp97

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 0.973001 mW
** Area: 6440 (mu_m)^2
** Transit frequency: 2.93601 MHz
** Transit frequency with error factor: 2.93561 MHz
** Slew rate: 3.80653 V/mu_s
** Phase margin: 88.8085°
** CMRR: 149 dB
** negPSRR: 49 dB
** posPSRR: 63 dB
** VoutMax: 4 V
** VoutMin: 0.370001 V
** VcmMax: 4.04001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -2.97409e+07 muA
** NormalTransistorNmos: 3.43181e+07 muA
** NormalTransistorNmos: 3.43171e+07 muA
** NormalTransistorNmos: 3.43181e+07 muA
** NormalTransistorNmos: 3.43171e+07 muA
** NormalTransistorPmos: -6.86369e+07 muA
** NormalTransistorPmos: -3.43189e+07 muA
** NormalTransistorPmos: -3.43189e+07 muA
** NormalTransistorNmos: 3.80921e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorPmos: -3.80929e+07 muA
** DiodeTransistorPmos: -3.80939e+07 muA
** NormalTransistorPmos: -3.80949e+07 muA
** NormalTransistorNmos: 3.80941e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** DiodeTransistorNmos: 2.97401e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24101  V
** in1: 2.5  V
** in2: 2.5  V
** inSourceTransconductanceComplementarySecondStage: 0.555001  V
** inStageBiasComplementarySecondStage: 4.21501  V
** innerComplementarySecondStage: 3.44001  V
** out: 2.5  V
** out1FirstStage: 0.555001  V
** out2FirstStage: 0.778001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 0.185001  V
** innerTransistorStack2Load1: 0.185001  V
** sourceTransconductance: 3.27001  V
** innerTransconductance: 0.150001  V
** inner: 0.150001  V


.END