.suckt  two_stage_single_output_op_amp_174_2 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos
m3 inputVoltageBiasXXpXX3 ibias sourceNmos sourceNmos nmos
m4 inputVoltageBiasXXnXX1 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m5 FirstStageYinnerSourceLoad1 inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m6 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m7 outFirstStage inputVoltageBiasXXpXX2 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m8 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos
m9 FirstStageYinnerSourceLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m10 FirstStageYinnerTransistorStack1Load2 ibias sourceNmos sourceNmos nmos
m11 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m12 FirstStageYinnerTransistorStack2Load2 ibias sourceNmos sourceNmos nmos
m13 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos
m14 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m15 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m16 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c2 out sourceNmos 
m17 out inputVoltageBiasXXnXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m18 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos
m19 out inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
m20 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m21 ibias ibias sourceNmos sourceNmos nmos
m22 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos
m23 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m24 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos
m25 inputVoltageBiasXXpXX3 inputVoltageBiasXXpXX3 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_174_2

