** Name: two_stage_single_output_op_amp_79_5

.MACRO two_stage_single_output_op_amp_79_5 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=36e-6
m2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=7e-6 W=51e-6
m3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=10e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=10e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=271e-6
m6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=108e-6
m7 inputVoltageBiasXXpXX2 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=231e-6
m8 out outFirstStage sourceNmos sourceNmos nmos4 L=1e-6 W=55e-6
m9 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=7e-6 W=339e-6
m10 outInputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=7e-6 W=53e-6
m11 FirstStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=7e-6 W=387e-6
m12 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=48e-6
m13 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=48e-6
m14 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=7e-6 W=339e-6
m15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=25e-6
m16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=25e-6
m17 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=7e-6 W=388e-6
m18 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=271e-6
m19 outFirstStage inputVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=144e-6
m20 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=262e-6
m21 FirstStageYout1 inputVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=144e-6
m22 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=249e-6
m23 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=249e-6
m24 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 8.30001e-12
.EOM two_stage_single_output_op_amp_79_5

** Expected Performance Values: 
** Gain: 127 dB
** Power consumption: 4.67901 mW
** Area: 14997 (mu_m)^2
** Transit frequency: 4.75201 MHz
** Transit frequency with error factor: 4.75218 MHz
** Slew rate: 10.8973 V/mu_s
** Phase margin: 60.1606°
** CMRR: 138 dB
** VoutMax: 3.86001 V
** VoutMin: 0.300001 V
** VcmMax: 5.22001 V
** VcmMin: 1.53001 V


** Expected Currents: 
** NormalTransistorNmos: 1.46741e+07 muA
** NormalTransistorNmos: 6.38641e+07 muA
** NormalTransistorPmos: -1.53269e+08 muA
** NormalTransistorPmos: -9.22399e+07 muA
** NormalTransistorPmos: -1.45065e+08 muA
** NormalTransistorPmos: -9.22399e+07 muA
** NormalTransistorPmos: -1.45065e+08 muA
** NormalTransistorNmos: 9.22391e+07 muA
** NormalTransistorNmos: 9.22381e+07 muA
** NormalTransistorNmos: 9.22391e+07 muA
** NormalTransistorNmos: 9.22381e+07 muA
** NormalTransistorNmos: 1.05651e+08 muA
** NormalTransistorNmos: 1.05652e+08 muA
** NormalTransistorNmos: 5.28251e+07 muA
** NormalTransistorNmos: 5.28251e+07 muA
** NormalTransistorNmos: 4.03881e+08 muA
** NormalTransistorPmos: -4.0388e+08 muA
** DiodeTransistorPmos: -4.03881e+08 muA
** DiodeTransistorNmos: 1.5327e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.46749e+07 muA
** NormalTransistorPmos: -1.46759e+07 muA
** DiodeTransistorPmos: -6.38649e+07 muA
** DiodeTransistorPmos: -6.38659e+07 muA


** Expected Voltages: 
** ibias: 0.556001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 3.09101  V
** out: 2.5  V
** outFirstStage: 0.701001  V
** outInputVoltageBiasXXpXX1: 3.29401  V
** outSourceVoltageBiasXXpXX1: 4.14801  V
** outSourceVoltageBiasXXpXX2: 4.25501  V
** outVoltageBiasXXnXX1: 0.906001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.351001  V
** innerTransistorStack1Load2: 0.351001  V
** innerTransistorStack2Load2: 0.351001  V
** out1: 0.555001  V
** sourceGCC1: 3.84401  V
** sourceGCC2: 3.84401  V
** sourceTransconductance: 1.67501  V
** inner: 4.14401  V


.END