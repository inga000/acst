** Name: two_stage_single_output_op_amp_38_10

.MACRO two_stage_single_output_op_amp_38_10 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=6e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=482e-6
mSimpleFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=50e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=26e-6
mMainBias5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
mSimpleFirstStageTransconductor6 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=16e-6
mSimpleFirstStageStageBias7 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=50e-6
mMainBias8 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=482e-6
mSecondStage1StageBias9 out ibias sourceNmos sourceNmos nmos4 L=3e-6 W=470e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=16e-6
mMainBias11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
mMainBias12 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=27e-6
mSimpleFirstStageLoad13 FirstStageYinnerSourceLoad1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=63e-6
mSimpleFirstStageLoad14 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=57e-6
mSimpleFirstStageLoad15 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=9e-6 W=57e-6
mSecondStage1Transconductor16 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=312e-6
mSecondStage1Transconductor17 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=600e-6
mSimpleFirstStageLoad18 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=63e-6
mMainBias19 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=10e-6 W=599e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 11.5e-12
.EOM two_stage_single_output_op_amp_38_10

** Expected Performance Values: 
** Gain: 102 dB
** Power consumption: 7.45601 mW
** Area: 14900 (mu_m)^2
** Transit frequency: 5.61201 MHz
** Transit frequency with error factor: 5.60949 MHz
** Slew rate: 5.28939 V/mu_s
** Phase margin: 60.1606°
** CMRR: 99 dB
** negPSRR: 110 dB
** posPSRR: 100 dB
** VoutMax: 4.25 V
** VoutMin: 0.240001 V
** VcmMax: 4.89001 V
** VcmMin: 1.44001 V


** Expected Currents: 
** NormalTransistorNmos: 2.46381e+07 muA
** NormalTransistorNmos: 4.50671e+07 muA
** NormalTransistorPmos: -5.76884e+08 muA
** NormalTransistorPmos: -3.04759e+07 muA
** NormalTransistorPmos: -3.04769e+07 muA
** NormalTransistorPmos: -3.04759e+07 muA
** NormalTransistorPmos: -3.04769e+07 muA
** NormalTransistorNmos: 6.09491e+07 muA
** DiodeTransistorNmos: 6.09481e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 3.04751e+07 muA
** NormalTransistorNmos: 7.73738e+08 muA
** NormalTransistorPmos: -7.73737e+08 muA
** NormalTransistorPmos: -7.73738e+08 muA
** DiodeTransistorNmos: 5.76885e+08 muA
** NormalTransistorNmos: 5.76885e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.46389e+07 muA
** DiodeTransistorPmos: -4.50679e+07 muA


** Expected Voltages: 
** ibias: 0.647001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 4.06401  V
** outInputVoltageBiasXXnXX1: 1.28801  V
** outSourceVoltageBiasXXnXX1: 0.644001  V
** outVoltageBiasXXpXX0: 3.70501  V
** outVoltageBiasXXpXX1: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 3.91801  V
** innerTransistorStack1Load1: 4.48201  V
** innerTransistorStack2Load1: 4.48201  V
** sourceTransconductance: 1.94501  V
** innerTransconductance: 4.62801  V
** inner: 0.644001  V


.END