** Name: two_stage_single_output_op_amp_36_9

.MACRO two_stage_single_output_op_amp_36_9 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=7e-6 W=7e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=8e-6 W=17e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=38e-6
m4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=600e-6
m5 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=51e-6
m6 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 pmos4 L=1e-6 W=67e-6
m7 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=58e-6
m8 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=7e-6 W=600e-6
m9 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=17e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=70e-6
m11 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=70e-6
m12 FirstStageYsourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=8e-6 W=38e-6
m13 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=8e-6 W=17e-6
m14 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=7e-6 W=7e-6
m15 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=329e-6
m16 outFirstStage FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=1e-6 W=67e-6
m17 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=62e-6
m18 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourcePmos sourcePmos pmos4 L=1e-6 W=58e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 9.20001e-12
.EOM two_stage_single_output_op_amp_36_9

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 4.86301 mW
** Area: 11427 (mu_m)^2
** Transit frequency: 7.65601 MHz
** Transit frequency with error factor: 7.65164 MHz
** Slew rate: 7.21554 V/mu_s
** Phase margin: 60.1606°
** CMRR: 109 dB
** negPSRR: 107 dB
** posPSRR: 100 dB
** VoutMax: 4.62001 V
** VoutMin: 1.09001 V
** VcmMax: 3.93001 V
** VcmMin: 1.77001 V


** Expected Currents: 
** NormalTransistorNmos: 2.42881e+07 muA
** NormalTransistorPmos: -2.93589e+07 muA
** DiodeTransistorPmos: -3.33319e+07 muA
** DiodeTransistorPmos: -3.33329e+07 muA
** NormalTransistorPmos: -3.33319e+07 muA
** NormalTransistorPmos: -3.33329e+07 muA
** NormalTransistorNmos: 6.66611e+07 muA
** DiodeTransistorNmos: 6.66601e+07 muA
** NormalTransistorNmos: 3.33311e+07 muA
** NormalTransistorNmos: 3.33311e+07 muA
** NormalTransistorNmos: 8.42257e+08 muA
** DiodeTransistorNmos: 8.42256e+08 muA
** NormalTransistorPmos: -8.42256e+08 muA
** DiodeTransistorNmos: 2.93581e+07 muA
** NormalTransistorNmos: 2.93581e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -2.42889e+07 muA


** Expected Voltages: 
** ibias: 1.49101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.00401  V
** out: 2.5  V
** outFirstStage: 4.05601  V
** outInputVoltageBiasXXnXX1: 1.62201  V
** outSourceVoltageBiasXXnXX1: 0.811001  V
** outSourceVoltageBiasXXnXX2: 0.747001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerOutputLoad1: 3.52501  V
** innerSourceLoad1: 4.25601  V
** innerTransistorStack2Load1: 4.25601  V
** sourceTransconductance: 1.94501  V
** inner: 0.811001  V
** inner: 0.741001  V


.END