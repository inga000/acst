** Name: two_stage_single_output_op_amp_16_3

.MACRO two_stage_single_output_op_amp_16_3 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=15e-6
m2 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=58e-6
m3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=4e-6 W=50e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=502e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=61e-6
m6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
m7 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=58e-6
m8 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=139e-6
m9 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=248e-6
m10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=35e-6
m11 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=4e-6 W=595e-6
m12 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=5e-6
m13 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=35e-6
m14 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=61e-6
m15 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=4e-6 W=35e-6
m16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=502e-6
Capacitor1 outFirstStage out 4.5e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_16_3

** Expected Performance Values: 
** Gain: 96 dB
** Power consumption: 1.74901 mW
** Area: 6552 (mu_m)^2
** Transit frequency: 2.51501 MHz
** Transit frequency with error factor: 2.50733 MHz
** Slew rate: 3.60026 V/mu_s
** Phase margin: 63.5984°
** CMRR: 94 dB
** negPSRR: 96 dB
** posPSRR: 144 dB
** VoutMax: 3.5 V
** VoutMin: 0.150001 V
** VcmMax: 3.23001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorNmos: 2.03879e+08 muA
** NormalTransistorPmos: -1.25019e+07 muA
** DiodeTransistorNmos: 1.22751e+07 muA
** NormalTransistorNmos: 1.22751e+07 muA
** NormalTransistorPmos: -2.45529e+07 muA
** DiodeTransistorPmos: -2.45539e+07 muA
** NormalTransistorPmos: -1.22759e+07 muA
** NormalTransistorPmos: -1.22759e+07 muA
** NormalTransistorNmos: 8.88421e+07 muA
** NormalTransistorPmos: -8.88429e+07 muA
** NormalTransistorPmos: -8.88419e+07 muA
** DiodeTransistorNmos: 1.25011e+07 muA
** DiodeTransistorPmos: -2.03878e+08 muA
** NormalTransistorPmos: -2.03879e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 2.91001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outInputVoltageBiasXXpXX1: 3.57201  V
** outSourceVoltageBiasXXpXX1: 4.28601  V
** outSourceVoltageBiasXXpXX2: 3.68601  V
** outVoltageBiasXXnXX0: 0.576001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** out1: 0.555001  V
** sourceTransconductance: 3.40601  V
** innerStageBias: 3.65601  V
** inner: 4.28601  V


.END