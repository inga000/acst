** Name: one_stage_single_output_op_amp89

.MACRO one_stage_single_output_op_amp89 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=9e-6
mMainBias3 ibias ibias sourcePmos sourcePmos pmos4 L=4e-6 W=36e-6
mMainBias4 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=8e-6 W=11e-6
mTelescopicFirstStageLoad5 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=107e-6
mTelescopicFirstStageLoad6 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=3e-6 W=107e-6
mTelescopicFirstStageLoad7 FirstStageYout1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=2e-6 W=71e-6
mTelescopicFirstStageLoad8 out inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=2e-6 W=71e-6
mMainBias9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=8e-6 W=17e-6
mTelescopicFirstStageLoad10 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=8e-6 W=95e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=296e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=2e-6 W=296e-6
mMainBias13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=68e-6
mTelescopicFirstStageLoad14 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=8e-6 W=95e-6
mMainBias15 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=4e-6 W=24e-6
mTelescopicFirstStageStageBias16 sourceTransconductance ibias sourcePmos sourcePmos pmos4 L=4e-6 W=528e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp89

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 0.974001 mW
** Area: 6560 (mu_m)^2
** Transit frequency: 6.73901 MHz
** Transit frequency with error factor: 6.73889 MHz
** Slew rate: 7.42969 V/mu_s
** Phase margin: 60.1606°
** CMRR: 145 dB
** VoutMax: 4.03001 V
** VoutMin: 0.300001 V
** VcmMax: 4.03001 V
** VcmMin: 0.150001 V


** Expected Currents: 
** NormalTransistorNmos: 1.27521e+07 muA
** NormalTransistorPmos: -6.76799e+06 muA
** NormalTransistorPmos: -1.91779e+07 muA
** NormalTransistorPmos: -6.80809e+07 muA
** NormalTransistorPmos: -6.80829e+07 muA
** NormalTransistorNmos: 6.80801e+07 muA
** NormalTransistorNmos: 6.80811e+07 muA
** NormalTransistorNmos: 6.80821e+07 muA
** NormalTransistorNmos: 6.80811e+07 muA
** NormalTransistorPmos: -1.48915e+08 muA
** NormalTransistorPmos: -6.80819e+07 muA
** NormalTransistorPmos: -6.80819e+07 muA
** DiodeTransistorNmos: 6.76701e+06 muA
** DiodeTransistorNmos: 1.91771e+07 muA
** DiodeTransistorPmos: -1.27529e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.18601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outVoltageBiasXXnXX0: 0.671001  V
** outVoltageBiasXXpXX1: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.22401  V
** innerTransistorStack1Load2: 0.150001  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.06401  V
** sourceGCC2: 3.06401  V


.END