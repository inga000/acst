** Name: two_stage_single_output_op_amp_114_12

.MACRO two_stage_single_output_op_amp_114_12 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos4 L=3e-6 W=7e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=146e-6
mTelescopicFirstStageStageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=173e-6
mSecondStage1StageBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=264e-6
mMainBias5 outVoltageBiasXXnXX3 outVoltageBiasXXnXX3 sourceTransconductance sourceTransconductance nmos4 L=5e-6 W=210e-6
mTelescopicFirstStageLoad6 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=7e-6 W=71e-6
mMainBias7 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=165e-6
mSecondStage1StageBias8 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=9e-6
mTelescopicFirstStageLoad9 FirstStageYout1 outVoltageBiasXXnXX3 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=5e-6 W=15e-6
mTelescopicFirstStageTransconductor10 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=9e-6
mTelescopicFirstStageTransconductor11 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=9e-6
mMainBias12 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=146e-6
mMainBias13 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias14 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=198e-6
mSecondStage1StageBias15 out ibias outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=3e-6 W=264e-6
mTelescopicFirstStageLoad16 outFirstStage outVoltageBiasXXnXX3 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=5e-6 W=15e-6
mMainBias17 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=3e-6 W=362e-6
mTelescopicFirstStageStageBias18 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=173e-6
mSecondStage1Transconductor19 SecondStageYinnerTransconductance outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=593e-6
mSecondStage1Transconductor20 out outVoltageBiasXXpXX1 SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=600e-6
mTelescopicFirstStageLoad21 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos4 L=7e-6 W=71e-6
mMainBias22 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=170e-6
mMainBias23 outVoltageBiasXXnXX3 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=192e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_114_12

** Expected Performance Values: 
** Gain: 149 dB
** Power consumption: 8.88001 mW
** Area: 9057 (mu_m)^2
** Transit frequency: 2.68101 MHz
** Transit frequency with error factor: 2.68027 MHz
** Slew rate: 14.9474 V/mu_s
** Phase margin: 74.4846°
** CMRR: 77 dB
** VoutMax: 4.55001 V
** VoutMin: 0.850001 V
** VcmMax: 4.51001 V
** VcmMin: 1.26001 V


** Expected Currents: 
** NormalTransistorNmos: 2.77914e+08 muA
** NormalTransistorNmos: 5.0767e+08 muA
** NormalTransistorPmos: -2.80885e+08 muA
** NormalTransistorPmos: -3.18072e+08 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** DiodeTransistorPmos: -5.71499e+06 muA
** NormalTransistorPmos: -5.71499e+06 muA
** NormalTransistorNmos: 3.29502e+08 muA
** DiodeTransistorNmos: 3.29502e+08 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 5.71401e+06 muA
** NormalTransistorNmos: 3.70071e+08 muA
** DiodeTransistorNmos: 3.70072e+08 muA
** NormalTransistorPmos: -3.7007e+08 muA
** NormalTransistorPmos: -3.70071e+08 muA
** DiodeTransistorNmos: 2.80886e+08 muA
** NormalTransistorNmos: 2.80885e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** NormalTransistorNmos: 9.99801e+06 muA
** DiodeTransistorNmos: 3.18073e+08 muA
** DiodeTransistorPmos: -2.77913e+08 muA
** DiodeTransistorPmos: -5.07669e+08 muA


** Expected Voltages: 
** ibias: 1.25601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX0: 4.00401  V
** out: 2.5  V
** outFirstStage: 4.24901  V
** outInputVoltageBiasXXnXX1: 1.11001  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXnXX2: 0.629001  V
** outVoltageBiasXXnXX3: 2.65001  V
** outVoltageBiasXXpXX1: 1.93601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** out1: 4.25801  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** innerTransconductance: 2.76201  V
** inner: 0.554001  V
** inner: 0.625  V


.END