** Name: symmetrical_op_amp37

.MACRO symmetrical_op_amp37 ibias in1 in2 out sourceNmos sourcePmos
m1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=17e-6
m2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
m3 inputVoltageBiasXXnXX0 inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=8e-6
m4 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
m5 ibias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=122e-6
m6 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
m7 inOutputStageBiasComplementarySecondStage inputVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=7e-6 W=43e-6
m8 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=6e-6 W=41e-6
m9 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=6e-6 W=41e-6
m10 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
m11 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=40e-6
m12 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=7e-6 W=512e-6
m13 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=28e-6
m14 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=2e-6 W=25e-6
m15 inputVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=7e-6 W=35e-6
m16 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=2e-6 W=31e-6
m17 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=2e-6 W=28e-6
m18 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=7e-6 W=272e-6
m19 FirstStageYsourceTransconductance inOutputStageBiasComplementarySecondStage FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=2e-6 W=15e-6
m20 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=98e-6
m21 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos4 L=2e-6 W=98e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp37

** Expected Performance Values: 
** Gain: 93 dB
** Power consumption: 0.863001 mW
** Area: 8512 (mu_m)^2
** Transit frequency: 2.59601 MHz
** Transit frequency with error factor: 2.596 MHz
** Slew rate: 3.5 V/mu_s
** Phase margin: 81.3601°
** CMRR: 144 dB
** negPSRR: 49 dB
** posPSRR: 58 dB
** VoutMax: 4.44001 V
** VoutMin: 0.420001 V
** VcmMax: 3.07001 V
** VcmMin: 0.0200001 V


** Expected Currents: 
** NormalTransistorNmos: 1.58251e+07 muA
** NormalTransistorPmos: -2.92399e+06 muA
** NormalTransistorPmos: -4.20899e+07 muA
** DiodeTransistorNmos: 1.12511e+07 muA
** DiodeTransistorNmos: 1.12491e+07 muA
** NormalTransistorPmos: -2.25009e+07 muA
** NormalTransistorPmos: -2.25019e+07 muA
** NormalTransistorPmos: -1.125e+07 muA
** NormalTransistorPmos: -1.125e+07 muA
** NormalTransistorNmos: 3.50261e+07 muA
** NormalTransistorNmos: 3.50251e+07 muA
** NormalTransistorPmos: -3.50269e+07 muA
** NormalTransistorPmos: -3.50259e+07 muA
** NormalTransistorPmos: -3.43319e+07 muA
** NormalTransistorPmos: -3.43329e+07 muA
** NormalTransistorNmos: 3.43311e+07 muA
** NormalTransistorNmos: 3.43301e+07 muA
** DiodeTransistorNmos: 2.92301e+06 muA
** DiodeTransistorNmos: 4.20891e+07 muA
** DiodeTransistorPmos: -1.58259e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25601  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 3.83801  V
** inOutputTransconductanceComplementarySecondStage: 0.826001  V
** inSourceTransconductanceComplementarySecondStage: 0.580001  V
** innerComplementarySecondStage: 4.23701  V
** inputVoltageBiasXXnXX0: 0.579001  V
** out: 2.5  V
** outFirstStage: 0.581001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 4.81001  V
** sourceTransconductance: 3.27501  V
** innerStageBias: 4.75901  V
** innerTransconductance: 0.176001  V
** inner: 4.79301  V
** inner: 0.177001  V


.END