.suckt  two_stage_fully_differential_op_amp_68_12 ibias in1 in2 out1 out2 sourceNmos sourcePmos vref
c_FullyDifferential_Compensation_Capacitor_1 out1FirstStage out1 
c_FullyDifferential_Compensation_Capacitor_2 out2FirstStage out2 
m_FullyDifferential_MainBias_1 inputVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX5 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_2 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX5 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_3 outInputVoltageBiasXXnXX1 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_4 outInputVoltageBiasXXnXX2 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_5 outInputVoltageBiasXXnXX3 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_6 outVoltageBiasXXnXX4 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_7 FeedbackStageYout1 FeedbackStageYout1 sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_Load_8 outFeedback outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FeedbackdStage_StageBias_9 FeedbackStageYsourceTransconductance1 ibias FeedbackStageYinnerStageBias1 FeedbackStageYinnerStageBias1 nmos
m_FullyDifferential_FeedbackdStage_StageBias_10 FeedbackStageYinnerStageBias1 outSourceVoltageBiasXXnXX5 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackdStage_StageBias_11 FeedbackStageYsourceTransconductance2 ibias FeedbackStageYinnerStageBias2 FeedbackStageYinnerStageBias2 nmos
m_FullyDifferential_FeedbackdStage_StageBias_12 FeedbackStageYinnerStageBias2 outSourceVoltageBiasXXnXX5 sourceNmos sourceNmos nmos
m_FullyDifferential_FeedbackStage_Transconductor_13 FeedbackStageYout1 out2 FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_14 outFeedback vref FeedbackStageYsourceTransconductance1 FeedbackStageYsourceTransconductance1 nmos
m_FullyDifferential_FeedbackStage_Transconductor_15 FeedbackStageYout1 out1 FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FeedbackStage_Transconductor_16 outFeedback vref FeedbackStageYsourceTransconductance2 FeedbackStageYsourceTransconductance2 nmos
m_FullyDifferential_FirstStage_Load_17 out1FirstStage outVoltageBiasXXnXX4 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m_FullyDifferential_FirstStage_Load_18 out2FirstStage outVoltageBiasXXnXX4 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m_FullyDifferential_FirstStage_Load_19 out1FirstStage outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_Load_20 out2FirstStage outFeedback sourcePmos sourcePmos pmos
m_FullyDifferential_FirstStage_StageBias_21 sourceTransconductance outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_FullyDifferential_FirstStage_StageBias_22 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_FirstStage_Transconductor_23 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m_FullyDifferential_FirstStage_Transconductor_24 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c_FullyDifferential_Load_Capacitor_3 out1 sourceNmos 
c_FullyDifferential_Load_Capacitor_4 out2 sourceNmos 
m_FullyDifferential_SecondStage1_StageBias_25 out1 outInputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos
m_FullyDifferential_SecondStage1_StageBias_26 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage1_Transconductor_27 out1 outVoltageBiasXXpXX1 SecondStage1YinnerTransconductance SecondStage1YinnerTransconductance pmos
m_FullyDifferential_SecondStage1_Transconductor_28 SecondStage1YinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage2_StageBias_29 out2 outInputVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos
m_FullyDifferential_SecondStage2_StageBias_30 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_SecondStage2_Transconductor_31 out2 outVoltageBiasXXpXX1 SecondStage2YinnerTransconductance SecondStage2YinnerTransconductance pmos
m_FullyDifferential_SecondStage2_Transconductor_32 SecondStage2YinnerTransconductance out2FirstStage sourcePmos sourcePmos pmos
m_FullyDifferential_MainBias_33 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos
m_FullyDifferential_MainBias_34 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_35 outInputVoltageBiasXXnXX2 outInputVoltageBiasXXnXX2 VoltageBiasXXnXX2Yinner VoltageBiasXXnXX2Yinner nmos
m_FullyDifferential_MainBias_36 VoltageBiasXXnXX2Yinner outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_37 outInputVoltageBiasXXnXX3 outInputVoltageBiasXXnXX3 VoltageBiasXXnXX3Yinner VoltageBiasXXnXX3Yinner nmos
m_FullyDifferential_MainBias_38 VoltageBiasXXnXX3Yinner outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_39 outVoltageBiasXXnXX4 outVoltageBiasXXnXX4 sourceTransconductance sourceTransconductance nmos
m_FullyDifferential_MainBias_40 ibias ibias outSourceVoltageBiasXXnXX5 outSourceVoltageBiasXXnXX5 nmos
m_FullyDifferential_MainBias_41 outSourceVoltageBiasXXnXX5 outSourceVoltageBiasXXnXX5 sourceNmos sourceNmos nmos
m_FullyDifferential_MainBias_42 inputVoltageBiasXXpXX0 inputVoltageBiasXXpXX0 sourcePmos sourcePmos pmos
m_FullyDifferential_SecondStage1_StageBias_43 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_fully_differential_op_amp_68_12

