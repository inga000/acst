** Name: two_stage_single_output_op_amp_44_8

.MACRO two_stage_single_output_op_amp_44_8 ibias in1 in2 out sourceNmos sourcePmos
m1 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=284e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=320e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=10e-6
m4 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=56e-6
m5 out outInputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=104e-6
m6 outFirstStage outInputVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=1e-6 W=10e-6
m7 FirstStageYout1 outInputVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=1e-6 W=10e-6
m8 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
m9 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=18e-6
m10 SecondStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=234e-6
m11 out outFirstStage sourcePmos sourcePmos pmos4 L=9e-6 W=398e-6
m12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=1e-6 W=19e-6
m13 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=599e-6
m14 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=4e-6 W=56e-6
m15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=29e-6
m16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=4e-6 W=29e-6
m17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=2e-6 W=24e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_44_8

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 5.73501 mW
** Area: 6545 (mu_m)^2
** Transit frequency: 2.81101 MHz
** Transit frequency with error factor: 2.81047 MHz
** Slew rate: 4.89342 V/mu_s
** Phase margin: 60.7336°
** CMRR: 136 dB
** VoutMax: 4.25 V
** VoutMin: 0.780001 V
** VcmMax: 3.79001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -6.0948e+08 muA
** NormalTransistorNmos: 2.20581e+07 muA
** NormalTransistorNmos: 3.42841e+07 muA
** NormalTransistorNmos: 2.20591e+07 muA
** NormalTransistorNmos: 3.42851e+07 muA
** NormalTransistorPmos: -2.20589e+07 muA
** NormalTransistorPmos: -2.20599e+07 muA
** DiodeTransistorPmos: -2.20589e+07 muA
** NormalTransistorPmos: -2.44529e+07 muA
** NormalTransistorPmos: -1.22269e+07 muA
** NormalTransistorPmos: -1.22269e+07 muA
** NormalTransistorNmos: 4.49006e+08 muA
** NormalTransistorNmos: 4.49005e+08 muA
** NormalTransistorPmos: -4.49005e+08 muA
** DiodeTransistorNmos: 6.09481e+08 muA
** DiodeTransistorNmos: 6.09482e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.10001  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.11901  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.14001  V
** out1: 3.32201  V
** sourceGCC1: 0.552001  V
** sourceGCC2: 0.552001  V
** sourceTransconductance: 3.37001  V
** innerStageBias: 0.488001  V


.END