** Name: two_stage_single_output_op_amp_101_3

.MACRO two_stage_single_output_op_amp_101_3 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=302e-6
m2 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=138e-6
m3 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=19e-6
m4 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=9e-6
m5 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
m6 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=216e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=237e-6
m8 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=2e-6 W=92e-6
m9 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=3e-6 W=138e-6
m10 out ibias SecondStageYinnerStageBias SecondStageYinnerStageBias pmos4 L=1e-6 W=565e-6
m11 outFirstStage inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=14e-6
m12 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=189e-6
m13 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=551e-6
m14 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=311e-6
m15 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=14e-6
m16 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=116e-6
m17 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=116e-6
m18 SecondStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=594e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 10.4001e-12
.EOM two_stage_single_output_op_amp_101_3

** Expected Performance Values: 
** Gain: 128 dB
** Power consumption: 5.62701 mW
** Area: 7823 (mu_m)^2
** Transit frequency: 5.80801 MHz
** Transit frequency with error factor: 5.80746 MHz
** Slew rate: 19.6977 V/mu_s
** Phase margin: 60.1606°
** CMRR: 128 dB
** VoutMax: 3.96001 V
** VoutMin: 0.300001 V
** VcmMax: 3 V
** VcmMin: 1.17001 V


** Expected Currents: 
** NormalTransistorNmos: 1.36363e+08 muA
** NormalTransistorPmos: -1.91622e+08 muA
** NormalTransistorPmos: -8.76139e+07 muA
** NormalTransistorPmos: -8.76139e+07 muA
** NormalTransistorNmos: 8.76131e+07 muA
** NormalTransistorNmos: 8.76131e+07 muA
** DiodeTransistorNmos: 8.76131e+07 muA
** NormalTransistorPmos: -3.11591e+08 muA
** NormalTransistorPmos: -3.11592e+08 muA
** NormalTransistorPmos: -8.76149e+07 muA
** NormalTransistorPmos: -8.76149e+07 muA
** NormalTransistorNmos: 6.02244e+08 muA
** NormalTransistorPmos: -6.02243e+08 muA
** NormalTransistorPmos: -6.02242e+08 muA
** DiodeTransistorNmos: 1.91623e+08 muA
** DiodeTransistorPmos: -1.36362e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.46301  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 1.36801  V
** out: 2.5  V
** outFirstStage: 0.705001  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.598001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.52201  V
** innerSourceLoad2: 0.555001  V
** innerStageBias: 4.20401  V
** out1: 1.11001  V
** sourceGCC1: 2.96201  V
** sourceGCC2: 2.95201  V
** innerStageBias: 4.27101  V


.END