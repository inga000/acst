** Name: two_stage_single_output_op_amp_48_9

.MACRO two_stage_single_output_op_amp_48_9 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 inputVoltageBiasXXnXX2 inputVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 nmos4 L=2e-6 W=34e-6
mMainBias2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=4e-6 W=10e-6
mSecondStage1StageBias3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=484e-6
mMainBias4 outSourceVoltageBiasXXnXX2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=40e-6
mFoldedCascodeFirstStageLoad5 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=84e-6
mFoldedCascodeFirstStageLoad6 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=4e-6 W=84e-6
mMainBias7 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=89e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 inputVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=13e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=30e-6
mMainBias11 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=10e-6
mSecondStage1StageBias12 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=484e-6
mFoldedCascodeFirstStageLoad13 outFirstStage inputVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=13e-6
mFoldedCascodeFirstStageLoad14 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=2e-6 W=84e-6
mFoldedCascodeFirstStageTransconductor15 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=106e-6
mFoldedCascodeFirstStageTransconductor16 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=6e-6 W=106e-6
mFoldedCascodeFirstStageStageBias17 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=6e-6 W=169e-6
mMainBias18 inputVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=335e-6
mSecondStage1Transconductor19 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=515e-6
mFoldedCascodeFirstStageLoad20 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=4e-6 W=84e-6
mMainBias21 outInputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=136e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_48_9

** Expected Performance Values: 
** Gain: 125 dB
** Power consumption: 4.39301 mW
** Area: 14531 (mu_m)^2
** Transit frequency: 3.88401 MHz
** Transit frequency with error factor: 3.88444 MHz
** Slew rate: 4.27068 V/mu_s
** Phase margin: 64.7443°
** CMRR: 142 dB
** VoutMax: 4.25 V
** VoutMin: 0.940001 V
** VcmMax: 4.07001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorPmos: -1.54699e+07 muA
** NormalTransistorPmos: -3.82219e+07 muA
** NormalTransistorNmos: 1.93331e+07 muA
** NormalTransistorNmos: 2.89981e+07 muA
** NormalTransistorNmos: 1.93351e+07 muA
** NormalTransistorNmos: 2.90001e+07 muA
** DiodeTransistorPmos: -1.93339e+07 muA
** NormalTransistorPmos: -1.93349e+07 muA
** NormalTransistorPmos: -1.93359e+07 muA
** DiodeTransistorPmos: -1.93349e+07 muA
** NormalTransistorPmos: -1.93319e+07 muA
** NormalTransistorPmos: -9.66599e+06 muA
** NormalTransistorPmos: -9.66599e+06 muA
** NormalTransistorNmos: 7.47e+08 muA
** DiodeTransistorNmos: 7.46999e+08 muA
** NormalTransistorPmos: -7.47e+08 muA
** DiodeTransistorNmos: 1.54691e+07 muA
** NormalTransistorNmos: 1.54681e+07 muA
** DiodeTransistorNmos: 3.82211e+07 muA
** DiodeTransistorNmos: 3.82201e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24101  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX2: 1.12401  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outInputVoltageBiasXXnXX1: 1.34801  V
** outSourceVoltageBiasXXnXX1: 0.674001  V
** outSourceVoltageBiasXXnXX2: 0.556001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.27501  V
** innerTransistorStack1Load2: 4.27301  V
** out1: 3.48301  V
** sourceGCC1: 0.531001  V
** sourceGCC2: 0.531001  V
** sourceTransconductance: 3.23901  V
** inner: 0.672001  V


.END