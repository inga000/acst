.suckt  two_stage_single_output_op_amp_93_1 ibias in1 in2 out sourceNmos sourcePmos
c_SingleOutput_Compensation_Capacitor_1 outFirstStage out 
m_SingleOutput_MainBias_1 outVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_2 outVoltageBiasXXnXX2 ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_3 FirstStageYout1 outVoltageBiasXXnXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos
m_SingleOutput_FirstStage_Load_4 outFirstStage outVoltageBiasXXnXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos
m_SingleOutput_FirstStage_Load_5 FirstStageYout1 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_6 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos
m_SingleOutput_FirstStage_Load_7 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_StageBias_8 sourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Transconductor_9 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos
m_SingleOutput_FirstStage_Transconductor_10 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos
c_SingleOutput_Load_Capacitor_2 out sourceNmos 
m_SingleOutput_SecondStage1_Transconductor_11 out outFirstStage sourceNmos sourceNmos nmos
m_SingleOutput_SecondStage1_StageBias_12 out ibias sourcePmos sourcePmos pmos
m_SingleOutput_MainBias_13 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceTransconductance sourceTransconductance nmos
m_SingleOutput_MainBias_14 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_15 ibias ibias sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_93_1

