** Name: two_stage_single_output_op_amp_99_1

.MACRO two_stage_single_output_op_amp_99_1 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=18e-6
m2 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=115e-6
m3 ibias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=31e-6
m4 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=52e-6
m5 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=3e-6 W=6e-6
m6 inputVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=190e-6
m7 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=513e-6
m8 outFirstStage FirstStageYout1 sourceNmos sourceNmos nmos4 L=8e-6 W=115e-6
m9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=5e-6 W=125e-6
m10 out ibias sourcePmos sourcePmos pmos4 L=2e-6 W=600e-6
m11 outFirstStage outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=4e-6
m12 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=2e-6 W=31e-6
m13 sourceTransconductance inputVoltageBiasXXpXX2 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=306e-6
m14 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=2e-6 W=394e-6
m15 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=4e-6
m16 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=136e-6
m17 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=136e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 11.6001e-12
.EOM two_stage_single_output_op_amp_99_1

** Expected Performance Values: 
** Gain: 100 dB
** Power consumption: 2.29601 mW
** Area: 9670 (mu_m)^2
** Transit frequency: 3.56201 MHz
** Transit frequency with error factor: 3.55903 MHz
** Slew rate: 6.13979 V/mu_s
** Phase margin: 60.1606°
** CMRR: 98 dB
** VoutMax: 4.81001 V
** VoutMin: 0.150001 V
** VcmMax: 3.32001 V
** VcmMin: 1.08001 V


** Expected Currents: 
** NormalTransistorNmos: 7.02521e+07 muA
** NormalTransistorNmos: 1.07627e+08 muA
** NormalTransistorPmos: -9.99599e+06 muA
** NormalTransistorPmos: -2.79339e+07 muA
** NormalTransistorPmos: -2.79339e+07 muA
** DiodeTransistorNmos: 2.79331e+07 muA
** NormalTransistorNmos: 2.79331e+07 muA
** NormalTransistorPmos: -1.26119e+08 muA
** NormalTransistorPmos: -1.2612e+08 muA
** NormalTransistorPmos: -2.79329e+07 muA
** NormalTransistorPmos: -2.79329e+07 muA
** NormalTransistorNmos: 1.95416e+08 muA
** NormalTransistorPmos: -1.95415e+08 muA
** DiodeTransistorNmos: 9.99501e+06 muA
** DiodeTransistorPmos: -7.02529e+07 muA
** DiodeTransistorPmos: -1.07626e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.24601  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.09401  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.587001  V
** outVoltageBiasXXpXX1: 1.31901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.27801  V
** innerStageBias: 4.81001  V
** out1: 0.556001  V
** sourceGCC1: 2.97101  V
** sourceGCC2: 2.97101  V


.END