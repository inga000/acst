** Name: two_stage_single_output_op_amp_12_8

.MACRO two_stage_single_output_op_amp_12_8 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=12e-6
mMainBias3 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=4e-6
mMainBias4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=435e-6
mSimpleFirstStageTransconductor5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=18e-6
mSimpleFirstStageStageBias6 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=3e-6 W=22e-6
mSecondStage1StageBias7 SecondStageYinnerStageBias ibias sourceNmos sourceNmos nmos4 L=3e-6 W=563e-6
mMainBias8 inputVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=13e-6
mSecondStage1StageBias9 out inputVoltageBiasXXnXX1 SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=1e-6 W=46e-6
mSimpleFirstStageTransconductor10 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=18e-6
mMainBias11 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=3e-6 W=272e-6
mSimpleFirstStageLoad12 FirstStageYinnerTransistorStack1Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=13e-6
mSimpleFirstStageLoad13 FirstStageYinnerTransistorStack2Load1 FirstStageYout1 sourcePmos sourcePmos pmos4 L=10e-6 W=13e-6
mSimpleFirstStageLoad14 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=4e-6 W=83e-6
mMainBias15 inputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=1e-6 W=523e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=146e-6
mSimpleFirstStageLoad17 outFirstStage inputVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=4e-6 W=83e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_12_8

** Expected Performance Values: 
** Gain: 91 dB
** Power consumption: 4.61701 mW
** Area: 5403 (mu_m)^2
** Transit frequency: 2.51001 MHz
** Transit frequency with error factor: 2.50796 MHz
** Slew rate: 3.69592 V/mu_s
** Phase margin: 64.7443°
** CMRR: 94 dB
** negPSRR: 95 dB
** posPSRR: 91 dB
** VoutMax: 4.30001 V
** VoutMin: 0.5 V
** VcmMax: 4.81001 V
** VcmMin: 0.800001 V


** Expected Currents: 
** NormalTransistorNmos: 2.08618e+08 muA
** NormalTransistorNmos: 1.00871e+07 muA
** NormalTransistorPmos: -2.47429e+08 muA
** NormalTransistorPmos: -8.36799e+06 muA
** NormalTransistorPmos: -8.36899e+06 muA
** NormalTransistorPmos: -8.36799e+06 muA
** NormalTransistorPmos: -8.36899e+06 muA
** NormalTransistorNmos: 1.67341e+07 muA
** NormalTransistorNmos: 8.36701e+06 muA
** NormalTransistorNmos: 8.36701e+06 muA
** NormalTransistorNmos: 4.30444e+08 muA
** NormalTransistorNmos: 4.30443e+08 muA
** NormalTransistorPmos: -4.30443e+08 muA
** DiodeTransistorNmos: 2.4743e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -2.08617e+08 muA
** DiodeTransistorPmos: -1.00879e+07 muA


** Expected Voltages: 
** ibias: 0.570001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.901001  V
** inputVoltageBiasXXpXX1: 3.68601  V
** out: 2.5  V
** outFirstStage: 3.73601  V
** outVoltageBiasXXpXX0: 4.27301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** out1: 3.83601  V
** sourceTransconductance: 1.86001  V
** innerStageBias: 0.165001  V


.END