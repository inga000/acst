** Name: symmetrical_op_amp116

.MACRO symmetrical_op_amp116 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias sourceNmos sourceNmos nmos4 L=10e-6 W=46e-6
m2 inOutputStageBiasComplementarySecondStage inOutputStageBiasComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=38e-6
m3 out2FirstStage out2FirstStage sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
m4 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=44e-6
m5 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=10e-6
m6 innerComplementarySecondStage inOutputStageBiasComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner nmos4 L=6e-6 W=22e-6
m7 out inOutputStageBiasComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias nmos4 L=6e-6 W=22e-6
m8 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=3e-6 W=10e-6
m9 out2FirstStage ibias sourceNmos sourceNmos nmos4 L=10e-6 W=116e-6
m10 outVoltageBiasXXpXX0 ibias sourceNmos sourceNmos nmos4 L=10e-6 W=56e-6
m11 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos4 L=10e-6 W=119e-6
m12 SecondStageYinnerStageBias innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=68e-6
m13 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourceNmos sourceNmos nmos4 L=6e-6 W=68e-6
m14 inOutputStageBiasComplementarySecondStage outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=2e-6 W=542e-6
m15 inSourceTransconductanceComplementarySecondStage out2FirstStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos4 L=2e-6 W=63e-6
m16 innerComplementarySecondStage out2FirstStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner pmos4 L=2e-6 W=174e-6
m17 out out2FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance pmos4 L=2e-6 W=174e-6
m18 out1FirstStage out2FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos4 L=2e-6 W=63e-6
m19 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=10e-6
m20 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=10e-6
m21 SecondStageYinnerTransconductance out1FirstStage sourcePmos sourcePmos pmos4 L=5e-6 W=27e-6
m22 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourcePmos sourcePmos pmos4 L=5e-6 W=27e-6
Capacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp116

** Expected Performance Values: 
** Gain: 95 dB
** Power consumption: 1.45501 mW
** Area: 7238 (mu_m)^2
** Transit frequency: 2.57401 MHz
** Transit frequency with error factor: 2.57369 MHz
** Slew rate: 3.50167 V/mu_s
** Phase margin: 82.506°
** CMRR: 138 dB
** negPSRR: 116 dB
** posPSRR: 62 dB
** VoutMax: 4.25 V
** VoutMin: 0.530001 V
** VcmMax: 4.81001 V
** VcmMin: 0.780001 V


** Expected Currents: 
** NormalTransistorNmos: 1.20161e+07 muA
** NormalTransistorNmos: 2.53821e+07 muA
** NormalTransistorPmos: -1.47983e+08 muA
** NormalTransistorPmos: -1.27669e+07 muA
** NormalTransistorPmos: -1.27679e+07 muA
** NormalTransistorPmos: -1.27669e+07 muA
** NormalTransistorPmos: -1.27679e+07 muA
** NormalTransistorNmos: 2.55331e+07 muA
** NormalTransistorNmos: 1.27661e+07 muA
** NormalTransistorNmos: 1.27661e+07 muA
** NormalTransistorNmos: 3.50901e+07 muA
** NormalTransistorNmos: 3.50891e+07 muA
** NormalTransistorPmos: -3.50909e+07 muA
** NormalTransistorPmos: -3.50899e+07 muA
** NormalTransistorNmos: 3.50901e+07 muA
** NormalTransistorNmos: 3.50891e+07 muA
** NormalTransistorPmos: -3.50909e+07 muA
** NormalTransistorPmos: -3.50899e+07 muA
** DiodeTransistorNmos: 1.47984e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorPmos: -1.20169e+07 muA
** DiodeTransistorPmos: -2.53829e+07 muA


** Expected Voltages: 
** ibias: 0.565001  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputStageBiasComplementarySecondStage: 0.931001  V
** inSourceTransconductanceComplementarySecondStage: 3.83601  V
** innerComplementarySecondStage: 0.596001  V
** out: 2.5  V
** out1FirstStage: 3.83601  V
** out2FirstStage: 3.68601  V
** outVoltageBiasXXpXX0: 4.26101  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load1: 4.40001  V
** innerTransistorStack2Load1: 4.40001  V
** sourceTransconductance: 1.88201  V
** innerStageBias: 0.191001  V
** innerTransconductance: 4.40001  V
** inner: 0.191001  V
** inner: 4.40001  V


.END