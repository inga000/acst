** Name: two_stage_single_output_op_amp_19_1

.MACRO two_stage_single_output_op_amp_19_1 ibias in1 in2 out sourceNmos sourcePmos
mSimpleFirstStageLoad1 FirstStageYinnerSourceLoad1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=49e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=25e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=4e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=50e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=13e-6
mSimpleFirstStageLoad6 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerSourceLoad1 sourceNmos sourceNmos nmos4 L=6e-6 W=49e-6
mMainBias7 inputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=92e-6
mSecondStage1Transconductor8 out outFirstStage sourceNmos sourceNmos nmos4 L=5e-6 W=297e-6
mSimpleFirstStageLoad9 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos4 L=10e-6 W=17e-6
mSimpleFirstStageTransconductor10 FirstStageYinnerSourceLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=19e-6
mSimpleFirstStageStageBias11 FirstStageYinnerStageBias ibias sourcePmos sourcePmos pmos4 L=3e-6 W=154e-6
mSimpleFirstStageStageBias12 FirstStageYsourceTransconductance inputVoltageBiasXXpXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=12e-6
mMainBias13 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=239e-6
mSecondStage1StageBias14 out ibias sourcePmos sourcePmos pmos4 L=3e-6 W=558e-6
mSimpleFirstStageTransconductor15 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=1e-6 W=19e-6
mMainBias16 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=3e-6 W=16e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 8.40001e-12
.EOM two_stage_single_output_op_amp_19_1

** Expected Performance Values: 
** Gain: 98 dB
** Power consumption: 1.45101 mW
** Area: 5895 (mu_m)^2
** Transit frequency: 2.75101 MHz
** Transit frequency with error factor: 2.7478 MHz
** Slew rate: 3.69939 V/mu_s
** Phase margin: 60.1606°
** CMRR: 103 dB
** negPSRR: 105 dB
** posPSRR: 156 dB
** VoutMax: 4.82001 V
** VoutMin: 0.150001 V
** VcmMax: 3.10001 V
** VcmMin: 0.320001 V


** Expected Currents: 
** NormalTransistorNmos: 7.42801e+07 muA
** NormalTransistorPmos: -3.25899e+06 muA
** NormalTransistorPmos: -4.78759e+07 muA
** DiodeTransistorNmos: 1.55551e+07 muA
** NormalTransistorNmos: 1.55551e+07 muA
** NormalTransistorNmos: 1.55551e+07 muA
** NormalTransistorPmos: -3.11129e+07 muA
** NormalTransistorPmos: -3.11139e+07 muA
** NormalTransistorPmos: -1.55559e+07 muA
** NormalTransistorPmos: -1.55559e+07 muA
** NormalTransistorNmos: 1.13667e+08 muA
** NormalTransistorPmos: -1.13666e+08 muA
** DiodeTransistorNmos: 3.25801e+06 muA
** DiodeTransistorNmos: 4.78751e+07 muA
** DiodeTransistorPmos: -7.42809e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.25201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.883001  V
** inputVoltageBiasXXpXX1: 3.86801  V
** out: 2.5  V
** outFirstStage: 0.555001  V
** outVoltageBiasXXnXX0: 0.575001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad1: 0.555001  V
** innerStageBias: 4.81101  V
** innerTransistorStack2Load1: 0.150001  V
** sourceTransconductance: 3.27701  V


.END