** Name: two_stage_single_output_op_amp_73_7

.MACRO two_stage_single_output_op_amp_73_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
mMainBias2 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=9e-6 W=11e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=37e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=3e-6 W=24e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=21e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=11e-6
mFoldedCascodeFirstStageLoad7 FirstStageYout1 FirstStageYinnerSourceLoad2 sourceNmos sourceNmos nmos4 L=6e-6 W=12e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=20e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=4e-6 W=20e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance outVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=9e-6 W=119e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=581e-6
mFoldedCascodeFirstStageLoad12 outFirstStage FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 nmos4 L=7e-6 W=67e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=3e-6 W=162e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=74e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=74e-6
mSecondStage1Transconductor16 out outFirstStage sourcePmos sourcePmos pmos4 L=1e-6 W=143e-6
mFoldedCascodeFirstStageLoad17 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=3e-6 W=162e-6
mMainBias18 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=123e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=3e-6 W=193e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.90001e-12
.EOM two_stage_single_output_op_amp_73_7

** Expected Performance Values: 
** Gain: 122 dB
** Power consumption: 8.47501 mW
** Area: 7730 (mu_m)^2
** Transit frequency: 4.93201 MHz
** Transit frequency with error factor: 4.93218 MHz
** Slew rate: 4.41787 V/mu_s
** Phase margin: 60.1606°
** CMRR: 146 dB
** VoutMax: 4.25 V
** VoutMin: 0.390001 V
** VcmMax: 5.12001 V
** VcmMin: 1.54001 V


** Expected Currents: 
** NormalTransistorPmos: -5.87849e+07 muA
** NormalTransistorPmos: -9.24099e+07 muA
** NormalTransistorPmos: -2.19309e+07 muA
** NormalTransistorPmos: -3.59109e+07 muA
** NormalTransistorPmos: -2.19309e+07 muA
** NormalTransistorPmos: -3.59109e+07 muA
** NormalTransistorNmos: 2.19301e+07 muA
** NormalTransistorNmos: 2.19301e+07 muA
** DiodeTransistorNmos: 2.19301e+07 muA
** NormalTransistorNmos: 2.79571e+07 muA
** NormalTransistorNmos: 2.79561e+07 muA
** NormalTransistorNmos: 1.39791e+07 muA
** NormalTransistorNmos: 1.39791e+07 muA
** NormalTransistorNmos: 1.45194e+09 muA
** NormalTransistorPmos: -1.45193e+09 muA
** DiodeTransistorNmos: 5.87841e+07 muA
** DiodeTransistorNmos: 9.24091e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32301  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.15201  V
** outVoltageBiasXXnXX1: 1.15501  V
** outVoltageBiasXXnXX2: 0.791001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 0.764001  V
** innerStageBias: 0.592001  V
** out1: 1.33301  V
** sourceGCC1: 4.03701  V
** sourceGCC2: 4.03701  V
** sourceTransconductance: 1.91301  V


.END