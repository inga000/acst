** Name: two_stage_single_output_op_amp_46_5

.MACRO two_stage_single_output_op_amp_46_5 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=10e-6 W=27e-6
m2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=52e-6
m3 inputVoltageBiasXXpXX2 inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=16e-6
m4 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=2e-6 W=5e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=244e-6
m6 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=105e-6
m7 FirstStageYout1 FirstStageYout1 FirstStageYinnerSourceLoad2 FirstStageYinnerSourceLoad2 pmos4 L=3e-6 W=145e-6
m8 inputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=13e-6
m9 out outFirstStage sourceNmos sourceNmos nmos4 L=2e-6 W=35e-6
m10 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=10e-6 W=52e-6
m11 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=50e-6
m12 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=10e-6 W=52e-6
m13 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=197e-6
m14 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=197e-6
m15 out outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=244e-6
m16 outFirstStage FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=145e-6
m17 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerSourceLoad2 sourcePmos sourcePmos pmos4 L=3e-6 W=105e-6
m18 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=51e-6
m19 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=8e-6 W=51e-6
m20 FirstStageYsourceTransconductance inputVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=5e-6 W=162e-6
m21 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=5e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.70001e-12
.EOM two_stage_single_output_op_amp_46_5

** Expected Performance Values: 
** Gain: 123 dB
** Power consumption: 2.77701 mW
** Area: 10672 (mu_m)^2
** Transit frequency: 2.54401 MHz
** Transit frequency with error factor: 2.54402 MHz
** Slew rate: 5.24589 V/mu_s
** Phase margin: 60.1606°
** CMRR: 137 dB
** VoutMax: 3.52001 V
** VoutMin: 0.560001 V
** VcmMax: 3.90001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 9.52401e+06 muA
** NormalTransistorNmos: 2.50101e+06 muA
** NormalTransistorNmos: 2.48951e+07 muA
** NormalTransistorNmos: 3.75221e+07 muA
** NormalTransistorNmos: 2.48951e+07 muA
** NormalTransistorNmos: 3.75221e+07 muA
** DiodeTransistorPmos: -2.48959e+07 muA
** DiodeTransistorPmos: -2.48969e+07 muA
** NormalTransistorPmos: -2.48959e+07 muA
** NormalTransistorPmos: -2.48969e+07 muA
** NormalTransistorPmos: -2.52569e+07 muA
** NormalTransistorPmos: -1.26279e+07 muA
** NormalTransistorPmos: -1.26279e+07 muA
** NormalTransistorNmos: 4.5832e+08 muA
** NormalTransistorPmos: -4.58319e+08 muA
** DiodeTransistorPmos: -4.5832e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -9.52499e+06 muA
** NormalTransistorPmos: -9.52599e+06 muA
** DiodeTransistorPmos: -2.50199e+06 muA


** Expected Voltages: 
** ibias: 1.16901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX2: 4.22701  V
** out: 2.5  V
** outFirstStage: 0.964001  V
** outInputVoltageBiasXXpXX1: 2.95201  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 3.97601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerSourceLoad2: 4.23601  V
** innerTransistorStack2Load2: 4.23501  V
** out1: 3.50201  V
** sourceGCC1: 0.525001  V
** sourceGCC2: 0.525001  V
** sourceTransconductance: 3.39601  V
** inner: 3.97601  V


.END