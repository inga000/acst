** Name: symmetrical_op_amp14

.MACRO symmetrical_op_amp14 ibias in1 in2 out sourceNmos sourcePmos
mSecondStage1StageBias1 inOutputTransconductanceComplementarySecondStage inOutputTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=4e-6 W=11e-6
mSymmetricalFirstStageLoad2 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=17e-6
mSymmetricalFirstStageLoad3 outFirstStage outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=17e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=1e-6 W=21e-6
mSecondStage1StageBias5 inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias6 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos4 L=1e-6 W=17e-6
mSecondStage1Transconductor7 SecondStageYinnerTransconductance outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=52e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor8 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos4 L=3e-6 W=52e-6
mSecondStageWithVoltageBiasAsStageBiasTransconductor9 innerComplementarySecondStage inOutputTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos4 L=4e-6 W=16e-6
mSecondStage1Transconductor10 out inOutputTransconductanceComplementarySecondStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos4 L=4e-6 W=16e-6
mSymmetricalFirstStageStageBias11 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos4 L=1e-6 W=47e-6
mSecondStageWithVoltageBiasAsStageBiasStageBias12 StageBiasComplementarySecondStageYinner inSourceStageBiasComplementarySecondStage sourcePmos sourcePmos pmos4 L=1e-6 W=17e-6
mMainBias13 inOutputTransconductanceComplementarySecondStage ibias sourcePmos sourcePmos pmos4 L=1e-6 W=108e-6
mSymmetricalFirstStageTransconductor14 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=104e-6
mSecondStage1StageBias15 out innerComplementarySecondStage inSourceStageBiasComplementarySecondStage inSourceStageBiasComplementarySecondStage pmos4 L=1e-6 W=17e-6
mSymmetricalFirstStageTransconductor16 outFirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=5e-6 W=104e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM symmetrical_op_amp14

** Expected Performance Values: 
** Gain: 94 dB
** Power consumption: 0.827001 mW
** Area: 1870 (mu_m)^2
** Transit frequency: 3.16901 MHz
** Transit frequency with error factor: 3.16894 MHz
** Slew rate: 3.50001 V/mu_s
** Phase margin: 81.3601°
** CMRR: 147 dB
** negPSRR: 47 dB
** posPSRR: 51 dB
** VoutMax: 3.75 V
** VoutMin: 0.470001 V
** VcmMax: 4.10001 V
** VcmMin: -0.00999999 V


** Expected Currents: 
** NormalTransistorPmos: -5.24319e+07 muA
** DiodeTransistorNmos: 1.14071e+07 muA
** DiodeTransistorNmos: 1.14071e+07 muA
** NormalTransistorPmos: -2.28169e+07 muA
** NormalTransistorPmos: -1.14079e+07 muA
** NormalTransistorPmos: -1.14079e+07 muA
** NormalTransistorNmos: 3.50121e+07 muA
** NormalTransistorNmos: 3.50111e+07 muA
** NormalTransistorPmos: -3.50129e+07 muA
** DiodeTransistorPmos: -3.50139e+07 muA
** DiodeTransistorPmos: -3.51509e+07 muA
** NormalTransistorPmos: -3.51519e+07 muA
** NormalTransistorNmos: 3.51501e+07 muA
** NormalTransistorNmos: 3.51491e+07 muA
** DiodeTransistorNmos: 5.24311e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.27201  V
** in1: 2.5  V
** in2: 2.5  V
** inOutputTransconductanceComplementarySecondStage: 0.880001  V
** inSourceStageBiasComplementarySecondStage: 4.09501  V
** inSourceTransconductanceComplementarySecondStage: 0.559001  V
** innerComplementarySecondStage: 3.19001  V
** out: 2.5  V
** outFirstStage: 0.559001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.23901  V
** innerTransconductance: 0.154001  V
** inner: 4.09301  V
** inner: 0.154001  V


.END