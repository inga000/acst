.suckt  one_stage_single_output_op_amp140 ibias in1 in2 out sourceNmos sourcePmos
m_SingleOutput_MainBias_1 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_2 FirstStageYinnerOutputLoad1 FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 pmos
m_SingleOutput_FirstStage_Load_3 FirstStageYinnerTransistorStack1Load1 FirstStageYinnerOutputLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_4 out FirstStageYinnerOutputLoad1 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 pmos
m_SingleOutput_FirstStage_Load_5 FirstStageYinnerTransistorStack2Load1 FirstStageYinnerOutputLoad1 sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Load_6 FirstStageYinnerOutputLoad1 inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos
m_SingleOutput_FirstStage_Load_7 FirstStageYinnerTransistorStack1Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_Load_8 out inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos
m_SingleOutput_FirstStage_Load_9 FirstStageYinnerTransistorStack2Load2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_FirstStage_StageBias_10 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m_SingleOutput_FirstStage_Transconductor_11 FirstStageYinnerOutputLoad1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m_SingleOutput_FirstStage_Transconductor_12 out in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c_SingleOutput_Load_Capacitor_1 out sourceNmos 
m_SingleOutput_MainBias_13 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos
m_SingleOutput_MainBias_14 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos
m_SingleOutput_MainBias_15 ibias ibias sourcePmos sourcePmos pmos
.end one_stage_single_output_op_amp140

