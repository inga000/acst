** Name: one_stage_single_output_op_amp103

.MACRO one_stage_single_output_op_amp103 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=123e-6
mMainBias2 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=61e-6
mMainBias3 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=28e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=1e-6 W=16e-6
mMainBias5 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mMainBias6 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourceTransconductance sourceTransconductance pmos4 L=4e-6 W=4e-6
mTelescopicFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=1e-6 W=123e-6
mTelescopicFirstStageLoad8 out outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=1e-6 W=123e-6
mMainBias9 outVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=3e-6 W=8e-6
mTelescopicFirstStageStageBias10 FirstStageYinnerStageBias outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=481e-6
mTelescopicFirstStageLoad11 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=600e-6
mTelescopicFirstStageTransconductor12 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=365e-6
mTelescopicFirstStageTransconductor13 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=365e-6
mTelescopicFirstStageLoad14 out outVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=600e-6
mMainBias15 outVoltageBiasXXnXX0 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=72e-6
mMainBias16 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=1e-6 W=209e-6
mTelescopicFirstStageStageBias17 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias pmos4 L=1e-6 W=593e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp103

** Expected Performance Values: 
** Gain: 89 dB
** Power consumption: 3.93001 mW
** Area: 10451 (mu_m)^2
** Transit frequency: 8.73801 MHz
** Transit frequency with error factor: 8.73826 MHz
** Slew rate: 23.8134 V/mu_s
** Phase margin: 70.4739°
** CMRR: 142 dB
** VoutMax: 3.27001 V
** VoutMin: 0.300001 V
** VcmMax: 3 V
** VcmMin: 0.440001 V


** Expected Currents: 
** NormalTransistorNmos: 9.53401e+06 muA
** NormalTransistorPmos: -7.29989e+07 muA
** NormalTransistorPmos: -2.11899e+08 muA
** NormalTransistorPmos: -2.35772e+08 muA
** NormalTransistorPmos: -2.35772e+08 muA
** DiodeTransistorNmos: 2.35773e+08 muA
** NormalTransistorNmos: 2.35773e+08 muA
** NormalTransistorNmos: 2.35773e+08 muA
** NormalTransistorPmos: -4.81077e+08 muA
** NormalTransistorPmos: -4.81078e+08 muA
** NormalTransistorPmos: -2.35771e+08 muA
** NormalTransistorPmos: -2.35771e+08 muA
** DiodeTransistorNmos: 7.29981e+07 muA
** DiodeTransistorNmos: 2.119e+08 muA
** DiodeTransistorPmos: -9.53499e+06 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.44801  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outSourceVoltageBiasXXpXX2: 4.19901  V
** outVoltageBiasXXnXX0: 0.610001  V
** outVoltageBiasXXnXX1: 0.705001  V
** outVoltageBiasXXpXX1: 2.18901  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.48701  V
** innerStageBias: 4.22401  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.04901  V
** sourceGCC2: 3.04901  V


.END