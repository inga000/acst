** Name: two_stage_single_output_op_amp_121_9

.MACRO two_stage_single_output_op_amp_121_9 ibias in1 in2 out sourceNmos sourcePmos
m1 ibias ibias outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 nmos4 L=4e-6 W=15e-6
m2 outInputVoltageBiasXXnXX1 outInputVoltageBiasXXnXX1 VoltageBiasXXnXX1Yinner VoltageBiasXXnXX1Yinner nmos4 L=1e-6 W=35e-6
m3 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=513e-6
m4 outSourceVoltageBiasXXnXX3 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
m5 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceTransconductance sourceTransconductance nmos4 L=4e-6 W=119e-6
m6 outVoltageBiasXXpXX0 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=43e-6
m7 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=24e-6
m8 outFirstStage outVoltageBiasXXnXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=4e-6 W=36e-6
m9 out outInputVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=1e-6 W=513e-6
m10 outVoltageBiasXXpXX0 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=73e-6
m11 outVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=563e-6
m12 sourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=194e-6
m13 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX3 sourceNmos sourceNmos nmos4 L=4e-6 W=541e-6
m14 FirstStageYout1 outVoltageBiasXXnXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=4e-6 W=36e-6
m15 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=27e-6
m16 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance nmos4 L=3e-6 W=27e-6
m17 VoltageBiasXXnXX1Yinner outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=1e-6 W=35e-6
m18 outFirstStage outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=1e-6 W=13e-6
m19 out outFirstStage sourcePmos sourcePmos pmos4 L=7e-6 W=225e-6
m20 outInputVoltageBiasXXnXX1 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=191e-6
m21 outVoltageBiasXXnXX2 outVoltageBiasXXpXX0 sourcePmos sourcePmos pmos4 L=7e-6 W=277e-6
m22 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=92e-6
m23 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=5e-6 W=92e-6
m24 FirstStageYout1 outVoltageBiasXXpXX1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=1e-6 W=13e-6
Capacitor1 outFirstStage out 12.3001e-12
Capacitor2 out sourceNmos 20e-12
.EOM two_stage_single_output_op_amp_121_9

** Expected Performance Values: 
** Gain: 129 dB
** Power consumption: 14.9961 mW
** Area: 13772 (mu_m)^2
** Transit frequency: 2.95301 MHz
** Transit frequency with error factor: 2.95319 MHz
** Slew rate: 21.0018 V/mu_s
** Phase margin: 60.1606°
** CMRR: 132 dB
** VoutMax: 3 V
** VoutMin: 0.860001 V
** VcmMax: 5.03001 V
** VcmMin: 1.36001 V


** Expected Currents: 
** NormalTransistorNmos: 3.50201e+07 muA
** NormalTransistorNmos: 2.68077e+08 muA
** NormalTransistorPmos: -1.52491e+08 muA
** NormalTransistorPmos: -2.24407e+08 muA
** NormalTransistorNmos: 1.71421e+07 muA
** NormalTransistorNmos: 1.71421e+07 muA
** NormalTransistorPmos: -1.71429e+07 muA
** NormalTransistorPmos: -1.71439e+07 muA
** NormalTransistorPmos: -1.71429e+07 muA
** NormalTransistorPmos: -1.71439e+07 muA
** NormalTransistorNmos: 2.58691e+08 muA
** NormalTransistorNmos: 2.5869e+08 muA
** NormalTransistorNmos: 1.71421e+07 muA
** NormalTransistorNmos: 1.71421e+07 muA
** NormalTransistorNmos: 2.27488e+09 muA
** DiodeTransistorNmos: 2.27488e+09 muA
** NormalTransistorPmos: -2.27487e+09 muA
** DiodeTransistorNmos: 1.52492e+08 muA
** NormalTransistorNmos: 1.52492e+08 muA
** DiodeTransistorNmos: 2.24408e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -3.50209e+07 muA
** DiodeTransistorPmos: -2.68076e+08 muA


** Expected Voltages: 
** ibias: 1.13701  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 2.43601  V
** outInputVoltageBiasXXnXX1: 1.26601  V
** outSourceVoltageBiasXXnXX1: 0.633001  V
** outSourceVoltageBiasXXnXX3: 0.555001  V
** outVoltageBiasXXnXX2: 2.65001  V
** outVoltageBiasXXpXX0: 3.87401  V
** outVoltageBiasXXpXX1: 3.64301  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 1.94501  V
** innerStageBias: 0.480001  V
** innerTransistorStack1Load2: 4.47801  V
** innerTransistorStack2Load2: 4.47801  V
** out1: 4.20701  V
** sourceGCC1: 2.09501  V
** sourceGCC2: 2.09501  V
** inner: 0.633001  V


.END