** Name: two_stage_single_output_op_amp_75_7

.MACRO two_stage_single_output_op_amp_75_7 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=7e-6
mMainBias3 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=5e-6
mMainBias4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=11e-6
mMainBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=10e-6
mFoldedCascodeFirstStageStageBias6 FirstStageYinnerStageBias outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
mFoldedCascodeFirstStageLoad7 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=14e-6
mFoldedCascodeFirstStageTransconductor8 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=64e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=10e-6 W=64e-6
mFoldedCascodeFirstStageStageBias10 FirstStageYsourceTransconductance inputVoltageBiasXXnXX1 FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=3e-6 W=56e-6
mSecondStage1StageBias11 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=2e-6 W=404e-6
mFoldedCascodeFirstStageLoad12 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=63e-6
mFoldedCascodeFirstStageLoad13 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=100e-6
mFoldedCascodeFirstStageLoad14 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=62e-6
mMainBias16 inputVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=91e-6
mSecondStage1Transconductor17 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=476e-6
mFoldedCascodeFirstStageLoad18 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=100e-6
mMainBias19 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=20e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_75_7

** Expected Performance Values: 
** Gain: 120 dB
** Power consumption: 9.33901 mW
** Area: 4438 (mu_m)^2
** Transit frequency: 7.69301 MHz
** Transit frequency with error factor: 7.69249 MHz
** Slew rate: 8.94038 V/mu_s
** Phase margin: 64.7443°
** CMRR: 141 dB
** VoutMax: 4.25 V
** VoutMin: 0.310001 V
** VcmMax: 5.17001 V
** VcmMin: 1.49001 V


** Expected Currents: 
** NormalTransistorPmos: -9.08929e+07 muA
** NormalTransistorPmos: -2.02769e+07 muA
** NormalTransistorPmos: -4.06129e+07 muA
** NormalTransistorPmos: -6.28599e+07 muA
** NormalTransistorPmos: -4.06129e+07 muA
** NormalTransistorPmos: -6.28599e+07 muA
** DiodeTransistorNmos: 4.06121e+07 muA
** NormalTransistorNmos: 4.06121e+07 muA
** NormalTransistorNmos: 4.06121e+07 muA
** NormalTransistorNmos: 4.44911e+07 muA
** NormalTransistorNmos: 4.44901e+07 muA
** NormalTransistorNmos: 2.22461e+07 muA
** NormalTransistorNmos: 2.22461e+07 muA
** NormalTransistorNmos: 1.61101e+09 muA
** NormalTransistorPmos: -1.611e+09 muA
** DiodeTransistorNmos: 9.08921e+07 muA
** DiodeTransistorNmos: 2.02761e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.40901  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 1.08001  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.19901  V
** outVoltageBiasXXnXX2: 0.713001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.508001  V
** innerTransistorStack2Load2: 0.524001  V
** out1: 0.666001  V
** sourceGCC1: 4.12301  V
** sourceGCC2: 4.12301  V
** sourceTransconductance: 1.89201  V


.END