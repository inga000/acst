** Name: two_stage_single_output_op_amp_66_5

.MACRO two_stage_single_output_op_amp_66_5 ibias in1 in2 out sourceNmos sourcePmos
mMainBias1 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=2e-6 W=10e-6
mMainBias2 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=10e-6
mMainBias3 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=8e-6 W=169e-6
mMainBias4 outInputVoltageBiasXXpXX2 outInputVoltageBiasXXpXX2 VoltageBiasXXpXX2Yinner VoltageBiasXXpXX2Yinner pmos4 L=3e-6 W=13e-6
mFoldedCascodeFirstStageStageBias5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=277e-6
mSecondStage1StageBias6 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=277e-6
mMainBias7 outVoltageBiasXXpXX3 outVoltageBiasXXpXX3 sourcePmos sourcePmos pmos4 L=3e-6 W=12e-6
mFoldedCascodeFirstStageLoad8 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 nmos4 L=2e-6 W=15e-6
mFoldedCascodeFirstStageLoad9 FirstStageYsourceGCC1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mFoldedCascodeFirstStageLoad10 FirstStageYsourceGCC2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=29e-6
mSecondStage1Transconductor11 out outFirstStage sourceNmos sourceNmos nmos4 L=3e-6 W=78e-6
mFoldedCascodeFirstStageLoad12 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 nmos4 L=2e-6 W=15e-6
mMainBias13 outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=12e-6
mMainBias14 outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=27e-6
mMainBias15 outVoltageBiasXXpXX3 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=2e-6 W=41e-6
mFoldedCascodeFirstStageLoad16 FirstStageYinnerTransistorStack1Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=67e-6
mFoldedCascodeFirstStageLoad17 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourcePmos sourcePmos pmos4 L=8e-6 W=67e-6
mFoldedCascodeFirstStageLoad18 FirstStageYout1 outVoltageBiasXXpXX3 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 pmos4 L=3e-6 W=83e-6
mFoldedCascodeFirstStageTransconductor19 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=175e-6
mFoldedCascodeFirstStageTransconductor20 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos4 L=10e-6 W=175e-6
mFoldedCascodeFirstStageStageBias21 FirstStageYsourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=8e-6 W=277e-6
mMainBias22 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=8e-6 W=169e-6
mMainBias23 VoltageBiasXXpXX2Yinner outSourceVoltageBiasXXpXX2 sourcePmos sourcePmos pmos4 L=3e-6 W=13e-6
mSecondStage1StageBias24 out outInputVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 outSourceVoltageBiasXXpXX2 pmos4 L=3e-6 W=277e-6
mFoldedCascodeFirstStageLoad25 outFirstStage outVoltageBiasXXpXX3 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 pmos4 L=3e-6 W=83e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_66_5

** Expected Performance Values: 
** Gain: 131 dB
** Power consumption: 3.51901 mW
** Area: 14592 (mu_m)^2
** Transit frequency: 3.86601 MHz
** Transit frequency with error factor: 3.86567 MHz
** Slew rate: 4.16226 V/mu_s
** Phase margin: 67.0361°
** CMRR: 139 dB
** VoutMax: 3.27001 V
** VoutMin: 0.510001 V
** VcmMax: 3.34001 V
** VcmMin: -0.409999 V


** Expected Currents: 
** NormalTransistorNmos: 1.17721e+07 muA
** NormalTransistorNmos: 2.64871e+07 muA
** NormalTransistorNmos: 4.06121e+07 muA
** NormalTransistorNmos: 1.88141e+07 muA
** NormalTransistorNmos: 2.84491e+07 muA
** NormalTransistorNmos: 1.88141e+07 muA
** NormalTransistorNmos: 2.84491e+07 muA
** NormalTransistorPmos: -1.88149e+07 muA
** NormalTransistorPmos: -1.88159e+07 muA
** NormalTransistorPmos: -1.88149e+07 muA
** NormalTransistorPmos: -1.88159e+07 muA
** NormalTransistorPmos: -1.92729e+07 muA
** DiodeTransistorPmos: -1.92739e+07 muA
** NormalTransistorPmos: -9.63599e+06 muA
** NormalTransistorPmos: -9.63599e+06 muA
** NormalTransistorNmos: 5.57932e+08 muA
** NormalTransistorPmos: -5.57931e+08 muA
** DiodeTransistorPmos: -5.57932e+08 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 9.99801e+06 muA
** DiodeTransistorPmos: -1.17729e+07 muA
** NormalTransistorPmos: -1.17739e+07 muA
** DiodeTransistorPmos: -2.64879e+07 muA
** NormalTransistorPmos: -2.64889e+07 muA
** DiodeTransistorPmos: -4.06129e+07 muA


** Expected Voltages: 
** ibias: 1.11601  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 0.911001  V
** outInputVoltageBiasXXpXX1: 3.51801  V
** outInputVoltageBiasXXpXX2: 2.70401  V
** outSourceVoltageBiasXXnXX1: 0.558001  V
** outSourceVoltageBiasXXpXX1: 4.25901  V
** outSourceVoltageBiasXXpXX2: 3.85201  V
** outVoltageBiasXXpXX3: 3.68601  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack1Load2: 4.44501  V
** innerTransistorStack2Load2: 4.44501  V
** out1: 4.08101  V
** sourceGCC1: 0.538001  V
** sourceGCC2: 0.538001  V
** sourceTransconductance: 3.23901  V
** inner: 4.25801  V
** inner: 3.85001  V


.END