** Name: one_stage_single_output_op_amp81

.MACRO one_stage_single_output_op_amp81 ibias in1 in2 out sourceNmos sourcePmos
mFoldedCascodeFirstStageLoad1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=41e-6
mFoldedCascodeFirstStageLoad2 FirstStageYout1 FirstStageYout1 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack1Load2 nmos4 L=10e-6 W=41e-6
mMainBias3 ibias ibias outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 nmos4 L=4e-6 W=4e-6
mMainBias4 outSourceVoltageBiasXXnXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=21e-6
mMainBias5 inputVoltageBiasXXpXX1 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=2e-6 W=5e-6
mMainBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=50e-6
mFoldedCascodeFirstStageStageBias7 FirstStageYinnerStageBias outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=160e-6
mFoldedCascodeFirstStageLoad8 FirstStageYinnerTransistorStack1Load2 FirstStageYinnerTransistorStack2Load2 sourceNmos sourceNmos nmos4 L=7e-6 W=41e-6
mFoldedCascodeFirstStageTransconductor9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageTransconductor10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=1e-6 W=20e-6
mFoldedCascodeFirstStageStageBias11 FirstStageYsourceTransconductance ibias FirstStageYinnerStageBias FirstStageYinnerStageBias nmos4 L=4e-6 W=34e-6
mMainBias12 inputVoltageBiasXXpXX1 outSourceVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=4e-6 W=38e-6
mFoldedCascodeFirstStageLoad13 out FirstStageYout1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=41e-6
mFoldedCascodeFirstStageLoad14 FirstStageYout1 inputVoltageBiasXXpXX1 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=2e-6 W=361e-6
mFoldedCascodeFirstStageLoad15 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=308e-6
mFoldedCascodeFirstStageLoad16 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=2e-6 W=308e-6
mFoldedCascodeFirstStageLoad17 out inputVoltageBiasXXpXX1 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=2e-6 W=361e-6
mLoadCapacitor1 out sourceNmos 20e-12
.EOM one_stage_single_output_op_amp81

** Expected Performance Values: 
** Gain: 86 dB
** Power consumption: 1.25501 mW
** Area: 5248 (mu_m)^2
** Transit frequency: 4.02201 MHz
** Transit frequency with error factor: 4.02217 MHz
** Slew rate: 3.64758 V/mu_s
** Phase margin: 84.7978°
** CMRR: 137 dB
** VoutMax: 4.08001 V
** VoutMin: 1.25 V
** VcmMax: 5.20001 V
** VcmMin: 1.44001 V


** Expected Currents: 
** NormalTransistorNmos: 1.81371e+07 muA
** NormalTransistorPmos: -7.33069e+07 muA
** NormalTransistorPmos: -1.114e+08 muA
** NormalTransistorPmos: -7.33069e+07 muA
** NormalTransistorPmos: -1.114e+08 muA
** DiodeTransistorNmos: 7.33061e+07 muA
** NormalTransistorNmos: 7.33051e+07 muA
** NormalTransistorNmos: 7.33061e+07 muA
** DiodeTransistorNmos: 7.33051e+07 muA
** NormalTransistorNmos: 7.61851e+07 muA
** NormalTransistorNmos: 7.61861e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** NormalTransistorNmos: 3.80931e+07 muA
** DiodeTransistorNmos: 9.99901e+06 muA
** DiodeTransistorNmos: 1.00001e+07 muA
** DiodeTransistorPmos: -1.81379e+07 muA
** DiodeTransistorPmos: -1.81389e+07 muA


** Expected Voltages: 
** ibias: 1.30201  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXpXX1: 3.03601  V
** out: 2.5  V
** outSourceVoltageBiasXXnXX1: 0.555001  V
** outSourceVoltageBiasXXpXX1: 4.23401  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerStageBias: 0.570001  V
** innerTransistorStack1Load2: 0.785001  V
** innerTransistorStack2Load2: 0.788001  V
** out1: 1.65101  V
** sourceGCC1: 3.75  V
** sourceGCC2: 3.75  V
** sourceTransconductance: 1.94501  V


.END