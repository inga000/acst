** Name: two_stage_single_output_op_amp_52_7

.MACRO two_stage_single_output_op_amp_52_7 ibias in1 in2 out sourceNmos sourcePmos
m1 outVoltageBiasXXnXX1 outVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=10e-6 W=69e-6
m2 outVoltageBiasXXnXX2 outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
m3 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
m4 ibias ibias outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=4e-6 W=37e-6
m5 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=24e-6
m6 out outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=342e-6
m7 outFirstStage outVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=10e-6 W=53e-6
m8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=2e-6 W=11e-6
m9 FirstStageYsourceGCC1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=22e-6
m10 FirstStageYsourceGCC2 in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos4 L=7e-6 W=22e-6
m11 FirstStageYsourceTransconductance outVoltageBiasXXnXX2 sourceNmos sourceNmos nmos4 L=5e-6 W=5e-6
m12 out outFirstStage sourcePmos sourcePmos pmos4 L=3e-6 W=359e-6
m13 outFirstStage ibias FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=4e-6 W=159e-6
m14 outVoltageBiasXXnXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=456e-6
m15 outVoltageBiasXXnXX2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=41e-6
m16 FirstStageYout1 ibias FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=4e-6 W=159e-6
m17 FirstStageYsourceGCC1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=59e-6
m18 FirstStageYsourceGCC2 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=4e-6 W=59e-6
Capacitor1 out sourceNmos 20e-12
Capacitor2 outFirstStage out 4.5e-12
.EOM two_stage_single_output_op_amp_52_7

** Expected Performance Values: 
** Gain: 121 dB
** Power consumption: 7.39101 mW
** Area: 8385 (mu_m)^2
** Transit frequency: 3.34401 MHz
** Transit frequency with error factor: 3.34352 MHz
** Slew rate: 3.54026 V/mu_s
** Phase margin: 61.3065°
** CMRR: 145 dB
** VoutMax: 4.25 V
** VoutMin: 0.450001 V
** VcmMax: 5.10001 V
** VcmMin: 1.04001 V


** Expected Currents: 
** NormalTransistorPmos: -1.91202e+08 muA
** NormalTransistorPmos: -1.71999e+07 muA
** NormalTransistorPmos: -1.61429e+07 muA
** NormalTransistorPmos: -2.47669e+07 muA
** NormalTransistorPmos: -1.61429e+07 muA
** NormalTransistorPmos: -2.47669e+07 muA
** DiodeTransistorNmos: 1.61421e+07 muA
** NormalTransistorNmos: 1.61421e+07 muA
** NormalTransistorNmos: 1.61421e+07 muA
** NormalTransistorNmos: 1.72451e+07 muA
** NormalTransistorNmos: 8.62301e+06 muA
** NormalTransistorNmos: 8.62301e+06 muA
** NormalTransistorNmos: 1.20018e+09 muA
** NormalTransistorPmos: -1.20017e+09 muA
** DiodeTransistorNmos: 1.91203e+08 muA
** DiodeTransistorNmos: 1.71991e+07 muA
** DiodeTransistorPmos: -9.99899e+06 muA
** DiodeTransistorPmos: -1e+07 muA


** Expected Voltages: 
** ibias: 3.32201  V
** in1: 2.5  V
** in2: 2.5  V
** out: 2.5  V
** outFirstStage: 3.68601  V
** outSourceVoltageBiasXXpXX1: 4.13101  V
** outVoltageBiasXXnXX1: 0.980001  V
** outVoltageBiasXXnXX2: 0.858001  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** innerTransistorStack2Load2: 0.386001  V
** out1: 0.591001  V
** sourceGCC1: 4.03601  V
** sourceGCC2: 4.03601  V
** sourceTransconductance: 1.91501  V


.END