.suckt  symmetrical_op_amp103 ibias in1 in2 out sourceNmos sourcePmos
m1 out1FirstStage out1FirstStage FirstStageYinnerTransistorStack1Load1 FirstStageYinnerTransistorStack1Load1 nmos
m2 FirstStageYinnerTransistorStack1Load1 out1FirstStage sourceNmos sourceNmos nmos
m3 inSourceTransconductanceComplementarySecondStage inSourceTransconductanceComplementarySecondStage FirstStageYinnerTransistorStack2Load1 FirstStageYinnerTransistorStack2Load1 nmos
m4 FirstStageYinnerTransistorStack2Load1 inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m5 FirstStageYsourceTransconductance ibias sourcePmos sourcePmos pmos
m6 out1FirstStage in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
m7 inSourceTransconductanceComplementarySecondStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance pmos
c1 out sourceNmos 
m8 out out1FirstStage SecondStageYinnerTransconductance SecondStageYinnerTransconductance nmos
m9 SecondStageYinnerTransconductance out1FirstStage sourceNmos sourceNmos nmos
m10 out innerComplementarySecondStage SecondStageYinnerStageBias SecondStageYinnerStageBias pmos
m11 SecondStageYinnerStageBias innerComplementarySecondStage sourcePmos sourcePmos pmos
m12 innerComplementarySecondStage innerComplementarySecondStage StageBiasComplementarySecondStageYinner StageBiasComplementarySecondStageYinner pmos
m13 StageBiasComplementarySecondStageYinner innerComplementarySecondStage sourcePmos sourcePmos pmos
m14 innerComplementarySecondStage inSourceTransconductanceComplementarySecondStage TransconductanceComplementarySecondStageYinner TransconductanceComplementarySecondStageYinner nmos
m15 TransconductanceComplementarySecondStageYinner inSourceTransconductanceComplementarySecondStage sourceNmos sourceNmos nmos
m16 ibias ibias sourcePmos sourcePmos pmos
.end symmetrical_op_amp103

