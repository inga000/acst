.suckt  two_stage_single_output_op_amp_8_1 ibias in1 in2 out sourceNmos sourcePmos
c1 outFirstStage out 
m1 outVoltageBiasXXpXX1 ibias sourceNmos sourceNmos nmos
m2 FirstStageYout1 FirstStageYout1 sourcePmos sourcePmos pmos
m3 outFirstStage FirstStageYout1 sourcePmos sourcePmos pmos
m4 FirstStageYsourceTransconductance ibias sourceNmos sourceNmos nmos
m5 FirstStageYout1 in1 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
m6 outFirstStage in2 FirstStageYsourceTransconductance FirstStageYsourceTransconductance nmos
c2 out sourceNmos 
m7 out outFirstStage sourceNmos sourceNmos nmos
m8 out outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
m9 ibias ibias sourceNmos sourceNmos nmos
m10 outVoltageBiasXXpXX1 outVoltageBiasXXpXX1 sourcePmos sourcePmos pmos
.end two_stage_single_output_op_amp_8_1

