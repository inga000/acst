** Name: two_stage_single_output_op_amp_104_1

.MACRO two_stage_single_output_op_amp_104_1 ibias in1 in2 out sourceNmos sourcePmos
mTelescopicFirstStageLoad1 FirstStageYout1 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=107e-6
mMainBias2 inputVoltageBiasXXnXX1 inputVoltageBiasXXnXX1 sourceNmos sourceNmos nmos4 L=3e-6 W=29e-6
mMainBias3 outVoltageBiasXXnXX0 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=56e-6
mMainBias4 ibias ibias sourcePmos sourcePmos pmos4 L=6e-6 W=36e-6
mMainBias5 outInputVoltageBiasXXpXX1 outInputVoltageBiasXXpXX1 VoltageBiasXXpXX1Yinner VoltageBiasXXpXX1Yinner pmos4 L=1e-6 W=43e-6
mTelescopicFirstStageStageBias6 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=436e-6
mMainBias7 outVoltageBiasXXpXX2 outVoltageBiasXXpXX2 sourceTransconductance sourceTransconductance pmos4 L=1e-6 W=14e-6
mTelescopicFirstStageLoad8 FirstStageYinnerTransistorStack2Load2 FirstStageYout1 sourceNmos sourceNmos nmos4 L=9e-6 W=107e-6
mSecondStage1Transconductor9 out outFirstStage sourceNmos sourceNmos nmos4 L=9e-6 W=393e-6
mTelescopicFirstStageLoad10 outFirstStage inputVoltageBiasXXnXX1 FirstStageYinnerTransistorStack2Load2 FirstStageYinnerTransistorStack2Load2 nmos4 L=3e-6 W=36e-6
mMainBias11 outInputVoltageBiasXXpXX1 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=53e-6
mMainBias12 outVoltageBiasXXpXX2 outVoltageBiasXXnXX0 sourceNmos sourceNmos nmos4 L=6e-6 W=409e-6
mTelescopicFirstStageLoad13 FirstStageYout1 outVoltageBiasXXpXX2 FirstStageYsourceGCC1 FirstStageYsourceGCC1 pmos4 L=1e-6 W=34e-6
mTelescopicFirstStageTransconductor14 FirstStageYsourceGCC1 in1 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=29e-6
mTelescopicFirstStageTransconductor15 FirstStageYsourceGCC2 in2 sourceTransconductance sourceTransconductance pmos4 L=5e-6 W=29e-6
mMainBias16 VoltageBiasXXpXX1Yinner outSourceVoltageBiasXXpXX1 sourcePmos sourcePmos pmos4 L=1e-6 W=43e-6
mMainBias17 inputVoltageBiasXXnXX1 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=259e-6
mSecondStage1StageBias18 out ibias sourcePmos sourcePmos pmos4 L=6e-6 W=374e-6
mTelescopicFirstStageLoad19 outFirstStage outVoltageBiasXXpXX2 FirstStageYsourceGCC2 FirstStageYsourceGCC2 pmos4 L=1e-6 W=34e-6
mMainBias20 outVoltageBiasXXnXX0 ibias sourcePmos sourcePmos pmos4 L=6e-6 W=65e-6
mTelescopicFirstStageStageBias21 sourceTransconductance outInputVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 outSourceVoltageBiasXXpXX1 pmos4 L=1e-6 W=436e-6
mLoadCapacitor1 out sourceNmos 20e-12
mCompensationCapacitor2 outFirstStage out 5.80001e-12
.EOM two_stage_single_output_op_amp_104_1

** Expected Performance Values: 
** Gain: 138 dB
** Power consumption: 2.05801 mW
** Area: 14500 (mu_m)^2
** Transit frequency: 2.66201 MHz
** Transit frequency with error factor: 2.6617 MHz
** Slew rate: 4.05864 V/mu_s
** Phase margin: 60.1606°
** CMRR: 132 dB
** VoutMax: 4.69001 V
** VoutMin: 0.170001 V
** VcmMax: 3.10001 V
** VcmMin: 0.340001 V


** Expected Currents: 
** NormalTransistorNmos: 1.73461e+07 muA
** NormalTransistorNmos: 1.32097e+08 muA
** NormalTransistorPmos: -1.81989e+07 muA
** NormalTransistorPmos: -7.29179e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** NormalTransistorPmos: -2.28569e+07 muA
** DiodeTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorNmos: 2.28561e+07 muA
** NormalTransistorPmos: -1.77813e+08 muA
** DiodeTransistorPmos: -1.77814e+08 muA
** NormalTransistorPmos: -2.28579e+07 muA
** NormalTransistorPmos: -2.28579e+07 muA
** NormalTransistorNmos: 1.05354e+08 muA
** NormalTransistorPmos: -1.05353e+08 muA
** DiodeTransistorNmos: 1.81981e+07 muA
** DiodeTransistorNmos: 7.29171e+07 muA
** DiodeTransistorPmos: -1.73469e+07 muA
** NormalTransistorPmos: -1.73479e+07 muA
** DiodeTransistorPmos: -1.32096e+08 muA
** DiodeTransistorPmos: -9.99899e+06 muA


** Expected Voltages: 
** ibias: 4.13001  V
** in1: 2.5  V
** in2: 2.5  V
** inputVoltageBiasXXnXX1: 0.705001  V
** out: 2.5  V
** outFirstStage: 0.573001  V
** outInputVoltageBiasXXpXX1: 3.57001  V
** outSourceVoltageBiasXXpXX1: 4.28501  V
** outVoltageBiasXXnXX0: 0.557001  V
** outVoltageBiasXXpXX2: 2.24501  V
** sourceNmos: 0  V
** sourcePmos: 5  V
** sourceTransconductance: 3.53201  V
** innerTransistorStack2Load2: 0.150001  V
** out1: 0.555001  V
** sourceGCC1: 3.00301  V
** sourceGCC2: 3.00301  V
** inner: 4.28401  V


.END